	-- Project Name: Voice Synthesizer
	
	library IEEE;
	use IEEE.STD_LOGIC_1164.ALL;
	use IEEE.STD_LOGIC_ARITH.ALL;
	use IEEE.STD_LOGIC_UNSIGNED.ALL;
	use IEEE.NUMERIC_STD.ALL;
	-- recuired libraries are used

entity Voice_Synthesizer is
		Port( CLK 	      : in 	STD_LOGIC;  --5 MHz
				B_ONE			: in  STD_LOGIC;	--first audio button
			 --B_ZERO		: in  STD_LOGIC;
				B_BES			: in  STD_LOGIC;	--second audio button
				DAC_CS  		: out STD_LOGIC;	--chip select pin of DAC
				DAC_CLR     : out STD_LOGIC;	--clear pin of DAC
				SPI_MOSI    : out STD_LOGIC;	--MOSI bit of SPI
				SPI_SCK     : out STD_LOGIC;	--SCK bit of SPI
				SPI_SS_B    : out STD_LOGIC;	--SS bit of SPI
				AMP_CS      : out STD_LOGIC;  
				AD_CONV     : out STD_LOGIC;
				SF_CE0      : out STD_LOGIC;
				FPGA_INIT_B : out STD_LOGIC);
end Voice_Synthesizer;
				
architecture Behavioral of Voice_Synthesizer is
				type One  is array (0 to 5403) of STD_LOGIC_VECTOR(15 downto 0);
				type Zero is array (0 to 4846) of STD_LOGIC_VECTOR(15 downto 0);
				type Bes  is array (0 to 4660) of STD_LOGIC_VECTOR(15 downto 0);
				signal One_voice : One :=(x"494E",x"464F",x"4953",x"4654",x"0E00",x"0000",x"4C61",x"7666",x"3538",x"2E37",x"362E",x"3130",x"3000",x"6461",x"7461",x"162A",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0100",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0200",x"0000",x"FDFF",x"FDFF",x"FFFF",x"FFFF",x"FCFF",x"FDFF",x"FEFF",x"0100",x"0000",x"FFFF",x"0400",x"FDFF",x"FBFF",x"FBFF",x"FEFF",x"FFFF",x"0100",x"FEFF",x"FFFF",x"FCFF",x"FCFF",x"FCFF",x"0000",x"0400",x"0600",x"0400",x"0100",x"0600",x"0200",x"FFFF",x"0000",x"FFFF",x"FEFF",x"0000",x"0000",x"0000",x"0000",x"FFFF",x"FDFF",x"FFFF",x"0200",x"0200",x"0200",x"0200",x"FFFF",x"0100",x"FFFF",x"0400",x"0400",x"0100",x"FEFF",x"FFFF",x"0000",x"0400",x"0600",x"0800",x"0200",x"FFFF",x"0100",x"FEFF",x"0100",x"FFFF",x"FDFF",x"FFFF",x"FEFF",x"FDFF",x"0000",x"0000",x"FDFF",x"FEFF",x"FBFF",x"F9FF",x"F6FF",x"FAFF",x"FBFF",x"FAFF",x"FEFF",x"0100",x"0600",x"0800",x"0800",x"0600",x"0700",x"0400",x"0100",x"0200",x"0000",x"0300",x"0200",x"0300",x"0100",x"FEFF",x"0000",x"0200",x"0200",x"0300",x"FEFF",x"FDFF",x"FDFF",x"0000",x"FFFF",x"FAFF",x"FEFF",x"FDFF",x"F9FF",x"FCFF",x"FBFF",x"FAFF",x"FCFF",x"FCFF",x"FDFF",x"0300",x"0800",x"0400",x"0000",x"0000",x"0400",x"0500",x"0500",x"0900",x"0800",x"0300",x"FFFF",x"FBFF",x"FBFF",x"FBFF",x"FEFF",x"FFFF",x"FEFF",x"0100",x"FFFF",x"0000",x"FFFF",x"FDFF",x"0000",x"FFFF",x"0000",x"0200",x"0400",x"0100",x"0000",x"FEFF",x"FEFF",x"FEFF",x"FFFF",x"0200",x"0700",x"0800",x"0600",x"0600",x"FEFF",x"0000",x"0100",x"FAFF",x"FBFF",x"FAFF",x"FBFF",x"F7FF",x"F4FF",x"FAFF",x"FCFF",x"FEFF",x"0200",x"0300",x"0500",x"0500",x"0A00",x"0800",x"0500",x"0300",x"0200",x"0500",x"0600",x"0600",x"0500",x"0100",x"0300",x"FFFF",x"FAFF",x"FAFF",x"F9FF",x"F9FF",x"FBFF",x"FEFF",x"FEFF",x"0000",x"0100",x"0400",x"0600",x"0300",x"FDFF",x"F9FF",x"FCFF",x"F7FF",x"F7FF",x"F8FF",x"FBFF",x"FDFF",x"0200",x"0200",x"0100",x"0100",x"0400",x"0700",x"0300",x"0100",x"0100",x"FFFF",x"FBFF",x"FFFF",x"0100",x"0500",x"0700",x"0300",x"0200",x"FFFF",x"FDFF",x"FFFF",x"0100",x"FFFF",x"FDFF",x"FEFF",x"0000",x"0300",x"0300",x"0100",x"FEFF",x"0100",x"0200",x"0200",x"0200",x"0200",x"0600",x"0100",x"0000",x"0000",x"FFFF",x"0200",x"0000",x"0200",x"0300",x"0600",x"FEFF",x"FEFF",x"0000",x"FCFF",x"0200",x"FFFF",x"FDFF",x"FFFF",x"0000",x"0300",x"0500",x"0200",x"FFFF",x"FCFF",x"F8FF",x"F9FF",x"F7FF",x"F8FF",x"FCFF",x"FEFF",x"0100",x"0100",x"0400",x"0300",x"0400",x"0300",x"0100",x"0300",x"0300",x"0300",x"0200",x"0300",x"0200",x"0000",x"0000",x"FFFF",x"FAFF",x"FDFF",x"FDFF",x"FDFF",x"FCFF",x"FEFF",x"FEFF",x"FCFF",x"FCFF",x"0000",x"0600",x"0900",x"0A00",x"0900",x"0A00",x"0500",x"0200",x"0300",x"0200",x"FEFF",x"FFFF",x"0000",x"FFFF",x"FFFF",x"FEFF",x"0200",x"0200",x"FEFF",x"0200",x"0400",x"0200",x"FFFF",x"0100",x"0100",x"FEFF",x"F8FF",x"F4FF",x"F5FF",x"F4FF",x"F7FF",x"F6FF",x"F8FF",x"FEFF",x"FDFF",x"FAFF",x"FDFF",x"FCFF",x"FBFF",x"0000",x"0300",x"0200",x"0300",x"0000",x"0400",x"0500",x"0300",x"0700",x"0600",x"0800",x"0800",x"0400",x"FFFF",x"F8FF",x"F8FF",x"FBFF",x"FCFF",x"FEFF",x"0000",x"0200",x"0000",x"0300",x"0400",x"0000",x"0500",x"0600",x"0100",x"FEFF",x"FBFF",x"FBFF",x"FBFF",x"FBFF",x"FFFF",x"0400",x"0800",x"0700",x"0500",x"0300",x"FFFF",x"FFFF",x"0500",x"0300",x"0900",x"0C00",x"0B00",x"0A00",x"0500",x"0100",x"FAFF",x"FBFF",x"FAFF",x"F6FF",x"F8FF",x"F8FF",x"F8FF",x"FCFF",x"FAFF",x"F7FF",x"F7FF",x"F7FF",x"FDFF",x"FFFF",x"FFFF",x"FFFF",x"F9FF",x"FAFF",x"FAFF",x"FAFF",x"FBFF",x"FEFF",x"0300",x"FDFF",x"0000",x"FEFF",x"FDFF",x"0500",x"0800",x"0A00",x"0A00",x"0500",x"0100",x"0400",x"0400",x"0000",x"0200",x"0400",x"0A00",x"0D00",x"0D00",x"0D00",x"1100",x"1100",x"1000",x"0B00",x"0900",x"0B00",x"0B00",x"0E00",x"0700",x"0300",x"0400",x"FFFF",x"FBFF",x"FDFF",x"FBFF",x"FAFF",x"F8FF",x"F6FF",x"F2FF",x"EFFF",x"F4FF",x"F2FF",x"EEFF",x"EEFF",x"F4FF",x"F7FF",x"F5FF",x"F9FF",x"FBFF",x"F6FF",x"F6FF",x"F7FF",x"F7FF",x"FAFF",x"FDFF",x"FEFF",x"FFFF",x"0100",x"FDFF",x"FAFF",x"FDFF",x"FFFF",x"0100",x"0400",x"0500",x"0600",x"0400",x"0300",x"0200",x"0000",x"0500",x"0300",x"0200",x"0400",x"0300",x"0400",x"0500",x"FEFF",x"FDFF",x"FCFF",x"FDFF",x"FFFF",x"0200",x"0600",x"0800",x"0900",x"0800",x"0B00",x"0800",x"0900",x"0D00",x"0E00",x"0D00",x"0B00",x"0600",x"FEFF",x"0200",x"0700",x"0700",x"0600",x"0900",x"0700",x"0100",x"FCFF",x"FDFF",x"F9FF",x"FAFF",x"FDFF",x"FCFF",x"FCFF",x"FEFF",x"F9FF",x"F5FF",x"FBFF",x"FBFF",x"FBFF",x"FAFF",x"FAFF",x"F7FF",x"F5FF",x"F6FF",x"F7FF",x"FAFF",x"FBFF",x"F7FF",x"FCFF",x"FCFF",x"FEFF",x"0000",x"FEFF",x"0200",x"0200",x"0300",x"0600",x"0700",x"0500",x"0500",x"0100",x"FEFF",x"0300",x"FEFF",x"FFFF",x"0300",x"0000",x"FFFF",x"FCFF",x"FEFF",x"FCFF",x"FBFF",x"F8FF",x"FBFF",x"F5FF",x"F7FF",x"FBFF",x"FCFF",x"0500",x"0700",x"0700",x"0800",x"0800",x"0800",x"0800",x"0A00",x"0400",x"0300",x"0600",x"0200",x"0500",x"0500",x"0300",x"FDFF",x"FBFF",x"FAFF",x"FAFF",x"F9FF",x"F7FF",x"F6FF",x"F7FF",x"F8FF",x"FCFF",x"0000",x"0200",x"0600",x"0900",x"1000",x"0F00",x"0E00",x"0C00",x"0900",x"0800",x"0600",x"0600",x"0300",x"0400",x"0500",x"0400",x"0400",x"0500",x"0600",x"0800",x"0600",x"0100",x"0200",x"FDFF",x"FAFF",x"FEFF",x"FFFF",x"FFFF",x"0000",x"0000",x"FDFF",x"FCFF",x"FFFF",x"FEFF",x"0000",x"FDFF",x"0200",x"0000",x"0200",x"0400",x"0100",x"FAFF",x"F0FF",x"ECFF",x"E8FF",x"E8FF",x"EFFF",x"F4FF",x"FBFF",x"FCFF",x"FAFF",x"FDFF",x"FEFF",x"FDFF",x"FCFF",x"FAFF",x"FBFF",x"FAFF",x"F9FF",x"FBFF",x"FBFF",x"FEFF",x"0600",x"0900",x"0900",x"0C00",x"1000",x"1100",x"0800",x"0A00",x"0B00",x"0900",x"0700",x"0700",x"0500",x"0500",x"0400",x"0000",x"0100",x"FCFF",x"F5FF",x"F4FF",x"FAFF",x"FEFF",x"0300",x"0500",x"0300",x"0200",x"FDFF",x"FDFF",x"FFFF",x"FCFF",x"FFFF",x"FCFF",x"FAFF",x"F8FF",x"F9FF",x"F6FF",x"F7FF",x"FCFF",x"0200",x"0600",x"0500",x"0800",x"0900",x"0900",x"0900",x"0900",x"0900",x"0B00",x"0500",x"0300",x"0300",x"0000",x"FDFF",x"0000",x"0600",x"0800",x"0600",x"0A00",x"0700",x"0100",x"F9FF",x"F9FF",x"FCFF",x"0000",x"0100",x"FEFF",x"FDFF",x"FDFF",x"FBFF",x"F7FF",x"F6FF",x"FBFF",x"FFFF",x"0400",x"0400",x"0400",x"0500",x"0500",x"0300",x"0300",x"0900",x"0B00",x"0500",x"0000",x"0000",x"FDFF",x"F7FF",x"F5FF",x"F5FF",x"F1FF",x"F1FF",x"F5FF",x"F3FF",x"F2FF",x"F6FF",x"FAFF",x"FDFF",x"FCFF",x"FDFF",x"0400",x"0300",x"FFFF",x"FFFF",x"FFFF",x"0100",x"0000",x"0400",x"0D00",x"0C00",x"0800",x"0300",x"0000",x"FDFF",x"FEFF",x"FEFF",x"FCFF",x"FFFF",x"0100",x"0300",x"0400",x"0300",x"0200",x"0300",x"0100",x"0100",x"0300",x"0600",x"0300",x"0100",x"0000",x"0000",x"0200",x"0100",x"0200",x"0400",x"0600",x"0500",x"0A00",x"0800",x"0600",x"0800",x"0400",x"0000",x"0200",x"FEFF",x"FCFF",x"0100",x"FDFF",x"F8FF",x"FAFF",x"FDFF",x"FBFF",x"0000",x"FEFF",x"FFFF",x"0100",x"0100",x"0000",x"FFFF",x"FFFF",x"FCFF",x"FCFF",x"FBFF",x"F9FF",x"F8FF",x"FEFF",x"0100",x"0300",x"0200",x"0200",x"0300",x"0500",x"0600",x"0300",x"FEFF",x"FDFF",x"FBFF",x"FAFF",x"F7FF",x"F7FF",x"FAFF",x"FCFF",x"FCFF",x"0000",x"0300",x"0100",x"0500",x"0400",x"0300",x"FFFF",x"F8FF",x"FAFF",x"0100",x"0200",x"FDFF",x"FCFF",x"FBFF",x"FBFF",x"FDFF",x"FFFF",x"0300",x"0A00",x"0800",x"0600",x"0300",x"0200",x"0400",x"0700",x"0500",x"0B00",x"0D00",x"0F00",x"0E00",x"0500",x"0000",x"FBFF",x"FBFF",x"F9FF",x"FAFF",x"FDFF",x"FBFF",x"F9FF",x"F6FF",x"FAFF",x"FFFF",x"0100",x"0400",x"0500",x"0300",x"0B00",x"0700",x"0300",x"0000",x"0200",x"0200",x"FFFF",x"FFFF",x"0100",x"FFFF",x"FDFF",x"FEFF",x"0500",x"0700",x"0500",x"0300",x"0200",x"FFFF",x"FDFF",x"FFFF",x"0000",x"FAFF",x"F9FF",x"FCFF",x"F8FF",x"F2FF",x"F2FF",x"F0FF",x"F6FF",x"FBFF",x"FFFF",x"FEFF",x"FAFF",x"FFFF",x"FEFF",x"0200",x"0300",x"0100",x"0300",x"FDFF",x"0000",x"0100",x"FFFF",x"FEFF",x"FAFF",x"F8FF",x"FBFF",x"FDFF",x"FBFF",x"F8FF",x"F6FF",x"F7FF",x"F8FF",x"FDFF",x"0100",x"0500",x"0500",x"0400",x"0700",x"0800",x"0A00",x"0900",x"0A00",x"0700",x"0200",x"0300",x"0300",x"0500",x"0300",x"0700",x"0600",x"0300",x"0500",x"0100",x"0100",x"0400",x"0700",x"0200",x"0000",x"FDFF",x"FFFF",x"FFFF",x"FDFF",x"0000",x"FDFF",x"0200",x"0400",x"0100",x"0100",x"0400",x"0400",x"0200",x"0400",x"0600",x"0400",x"0000",x"0100",x"0100",x"0200",x"0300",x"0500",x"0500",x"0400",x"0100",x"FFFF",x"FEFF",x"FBFF",x"FAFF",x"FCFF",x"FEFF",x"0500",x"0700",x"0300",x"0400",x"FFFF",x"FBFF",x"FAFF",x"FBFF",x"FEFF",x"0100",x"FDFF",x"FBFF",x"FEFF",x"FEFF",x"FAFF",x"FBFF",x"FAFF",x"F6FF",x"F7FF",x"F8FF",x"F5FF",x"F8FF",x"F9FF",x"FAFF",x"FDFF",x"FBFF",x"FEFF",x"0500",x"0A00",x"0A00",x"0800",x"0400",x"0000",x"0000",x"FBFF",x"F9FF",x"F8FF",x"F9FF",x"FCFF",x"0100",x"0500",x"0B00",x"0F00",x"0F00",x"0D00",x"0B00",x"0900",x"0500",x"FFFF",x"F8FF",x"F8FF",x"F6FF",x"F4FF",x"F1FF",x"F1FF",x"F7FF",x"F8FF",x"FEFF",x"0600",x"0700",x"0700",x"0500",x"0400",x"0100",x"0600",x"0900",x"0700",x"0900",x"0C00",x"0C00",x"0B00",x"0600",x"0200",x"0600",x"0500",x"0500",x"0500",x"0300",x"0200",x"0100",x"0100",x"FCFF",x"FBFF",x"0200",x"0500",x"0700",x"0900",x"0600",x"0100",x"FCFF",x"F5FF",x"F1FF",x"EEFF",x"F5FF",x"F5FF",x"FBFF",x"FDFF",x"FDFF",x"FCFF",x"FAFF",x"FCFF",x"FEFF",x"FFFF",x"FFFF",x"FCFF",x"F9FF",x"FAFF",x"FAFF",x"FEFF",x"0300",x"0200",x"0800",x"0400",x"0100",x"0100",x"FFFF",x"0100",x"0300",x"0100",x"FEFF",x"FEFF",x"FDFF",x"FEFF",x"FBFF",x"FDFF",x"0400",x"0900",x"0C00",x"0700",x"0100",x"FEFF",x"F7FF",x"F3FF",x"F5FF",x"F8FF",x"FFFF",x"0400",x"0700",x"0500",x"0100",x"0000",x"0400",x"0200",x"0600",x"0900",x"0600",x"FDFF",x"FAFF",x"FEFF",x"FDFF",x"0100",x"0300",x"0100",x"0300",x"0300",x"0300",x"0100",x"0200",x"0600",x"0600",x"0300",x"0000",x"0100",x"0100",x"FEFF",x"F9FF",x"FAFF",x"F9FF",x"F9FF",x"FCFF",x"FEFF",x"FEFF",x"FBFF",x"FAFF",x"FAFF",x"FBFF",x"FBFF",x"0000",x"0400",x"0500",x"0400",x"0200",x"0400",x"0300",x"0200",x"0100",x"0100",x"0000",x"FAFF",x"FBFF",x"FEFF",x"0400",x"0900",x"0900",x"0B00",x"0A00",x"0800",x"0600",x"0500",x"0000",x"FAFF",x"FDFF",x"0000",x"0300",x"0700",x"0900",x"0600",x"0400",x"0000",x"FCFF",x"FBFF",x"FFFF",x"FEFF",x"FDFF",x"0200",x"0400",x"0500",x"0000",x"0000",x"0200",x"0100",x"FDFF",x"0100",x"0200",x"FFFF",x"FFFF",x"FFFF",x"0000",x"0000",x"0200",x"0200",x"0300",x"0400",x"FFFF",x"FEFF",x"FEFF",x"FFFF",x"FFFF",x"FBFF",x"F7FF",x"F5FF",x"F3FF",x"F6FF",x"FBFF",x"FAFF",x"FAFF",x"F8FF",x"F7FF",x"F5FF",x"F5FF",x"F8FF",x"F6FF",x"F7FF",x"F8FF",x"F7FF",x"FBFF",x"F8FF",x"F7FF",x"FCFF",x"0400",x"0700",x"0C00",x"0B00",x"0A00",x"0B00",x"0700",x"0700",x"0700",x"0900",x"0600",x"0700",x"0400",x"FFFF",x"FFFF",x"FDFF",x"FEFF",x"FFFF",x"FEFF",x"FDFF",x"0300",x"0400",x"0000",x"0100",x"0500",x"0500",x"0800",x"0B00",x"0600",x"0100",x"0500",x"0700",x"0400",x"0500",x"0500",x"0600",x"0800",x"0300",x"0300",x"0300",x"0300",x"0200",x"0100",x"FFFF",x"FBFF",x"0000",x"0400",x"FEFF",x"FAFF",x"FAFF",x"F8FF",x"F5FF",x"F9FF",x"FCFF",x"0000",x"0300",x"0100",x"0000",x"FEFF",x"F8FF",x"FAFF",x"FBFF",x"FCFF",x"FEFF",x"FDFF",x"FEFF",x"0000",x"0500",x"0300",x"FDFF",x"FBFF",x"FCFF",x"FFFF",x"0200",x"0400",x"0300",x"0200",x"0500",x"0300",x"FEFF",x"FDFF",x"FBFF",x"FBFF",x"F7FF",x"F6FF",x"FAFF",x"FAFF",x"FCFF",x"FCFF",x"0000",x"FBFF",x"FAFF",x"FAFF",x"FAFF",x"F6FF",x"F1FF",x"F6FF",x"FAFF",x"F8FF",x"FAFF",x"FCFF",x"FBFF",x"FDFF",x"FEFF",x"0200",x"0300",x"0600",x"0E00",x"1300",x"1700",x"1600",x"1400",x"1500",x"1600",x"1600",x"1300",x"0B00",x"0900",x"0600",x"FDFF",x"FBFF",x"F9FF",x"F7FF",x"FEFF",x"FDFF",x"FDFF",x"0000",x"FFFF",x"FDFF",x"0400",x"0600",x"0200",x"0300",x"0100",x"0000",x"FDFF",x"FCFF",x"FFFF",x"FDFF",x"0200",x"0400",x"0200",x"0600",x"0700",x"0500",x"0000",x"FDFF",x"F6FF",x"F2FF",x"F7FF",x"F6FF",x"F8FF",x"F4FF",x"F7FF",x"FDFF",x"F9FF",x"F3FF",x"F5FF",x"F7FF",x"FCFF",x"FFFF",x"0400",x"0900",x"0400",x"0200",x"FFFF",x"FBFF",x"FCFF",x"F9FF",x"FAFF",x"FEFF",x"FBFF",x"FEFF",x"0100",x"0400",x"0800",x"0300",x"0100",x"0400",x"FEFF",x"FEFF",x"0200",x"0200",x"0400",x"0500",x"0800",x"0500",x"0500",x"0500",x"0100",x"0100",x"0300",x"0200",x"0000",x"FDFF",x"FAFF",x"F7FF",x"F9FF",x"FCFF",x"FCFF",x"FAFF",x"F8FF",x"FAFF",x"FBFF",x"FFFF",x"FDFF",x"0000",x"0800",x"0800",x"0700",x"0700",x"0600",x"0900",x"0600",x"0500",x"0200",x"FCFF",x"FDFF",x"FFFF",x"0100",x"0400",x"0400",x"0400",x"0800",x"FFFF",x"FCFF",x"FCFF",x"F7FF",x"FBFF",x"FDFF",x"0100",x"0900",x"0700",x"0400",x"0300",x"0300",x"0500",x"0800",x"0800",x"0400",x"0200",x"0400",x"0300",x"0000",x"FEFF",x"0500",x"0900",x"0A00",x"0800",x"0000",x"FDFF",x"FBFF",x"F5FF",x"EFFF",x"F0FF",x"EFFF",x"EAFF",x"F5FF",x"FAFF",x"FEFF",x"0800",x"0B00",x"0C00",x"0900",x"0900",x"0600",x"0000",x"FAFF",x"FAFF",x"F6FF",x"F4FF",x"F7FF",x"F9FF",x"FDFF",x"FEFF",x"FDFF",x"FDFF",x"F7FF",x"F8FF",x"FFFF",x"F5FF",x"F8FF",x"0000",x"FDFF",x"FFFF",x"0100",x"0300",x"0300",x"0300",x"0300",x"0200",x"0000",x"0400",x"0800",x"0900",x"0800",x"0400",x"0200",x"0000",x"0500",x"0400",x"FFFF",x"0000",x"0000",x"0500",x"0900",x"0300",x"0400",x"0200",x"FEFF",x"FEFF",x"F9FF",x"0100",x"0900",x"0B00",x"1100",x"1400",x"1000",x"0C00",x"0300",x"0300",x"FFFF",x"F9FF",x"FBFF",x"FAFF",x"FCFF",x"F6FF",x"F4FF",x"FAFF",x"FEFF",x"0400",x"0600",x"0800",x"0800",x"0600",x"0300",x"FFFF",x"FEFF",x"FAFF",x"F1FF",x"F1FF",x"F4FF",x"F5FF",x"F8FF",x"FDFF",x"0100",x"0500",x"0A00",x"0600",x"FEFF",x"F9FF",x"FAFF",x"FDFF",x"FAFF",x"0100",x"0300",x"0100",x"0500",x"0000",x"FFFF",x"0100",x"FCFF",x"FBFF",x"FCFF",x"FEFF",x"FFFF",x"FFFF",x"FFFF",x"0400",x"0800",x"0300",x"0100",x"FFFF",x"F8FF",x"F2FF",x"F5FF",x"F9FF",x"F9FF",x"FAFF",x"F8FF",x"FDFF",x"0400",x"0100",x"0300",x"0800",x"1100",x"1300",x"0E00",x"0D00",x"0B00",x"0900",x"0600",x"0000",x"0100",x"0200",x"0000",x"FFFF",x"FCFF",x"F6FF",x"F5FF",x"FEFF",x"FEFF",x"0100",x"0000",x"0300",x"FCFF",x"F9FF",x"F9FF",x"F9FF",x"FFFF",x"0600",x"0400",x"0700",x"0200",x"0300",x"0500",x"0000",x"FFFF",x"FEFF",x"F8FF",x"F2FF",x"F4FF",x"F5FF",x"FBFF",x"0100",x"0200",x"0500",x"0400",x"0200",x"0800",x"0700",x"FCFF",x"F9FF",x"F5FF",x"F4FF",x"F8FF",x"F9FF",x"0200",x"0600",x"0C00",x"0C00",x"0B00",x"0C00",x"0C00",x"0800",x"0300",x"0200",x"0000",x"FBFF",x"0100",x"0300",x"FFFF",x"0300",x"0500",x"0800",x"0600",x"0300",x"0300",x"0100",x"0000",x"FEFF",x"0200",x"0400",x"0400",x"0400",x"0400",x"0700",x"0900",x"0600",x"FFFF",x"FBFF",x"F8FF",x"F6FF",x"F4FF",x"EDFF",x"EEFF",x"F1FF",x"F1FF",x"F3FF",x"F8FF",x"F8FF",x"FBFF",x"FDFF",x"F9FF",x"0100",x"0300",x"0100",x"0200",x"FCFF",x"FCFF",x"F9FF",x"FAFF",x"0100",x"0100",x"0400",x"0400",x"0800",x"0600",x"FDFF",x"FCFF",x"FAFF",x"FEFF",x"0400",x"0600",x"0500",x"0000",x"0200",x"0600",x"0700",x"0600",x"0B00",x"0E00",x"1000",x"1100",x"0B00",x"0300",x"FFFF",x"FFFF",x"FEFF",x"FFFF",x"0400",x"0200",x"0100",x"0600",x"0500",x"0100",x"FCFF",x"F7FF",x"F7FF",x"F4FF",x"F2FF",x"F7FF",x"FAFF",x"FEFF",x"0300",x"FEFF",x"FCFF",x"0000",x"FEFF",x"F8FF",x"FAFF",x"FFFF",x"0200",x"0300",x"0700",x"0700",x"0400",x"0500",x"0300",x"0200",x"0300",x"0000",x"0300",x"FEFF",x"FAFF",x"FAFF",x"FBFF",x"FCFF",x"F7FF",x"F7FF",x"FDFF",x"FFFF",x"FDFF",x"0200",x"0200",x"0400",x"0500",x"0500",x"0900",x"0B00",x"0A00",x"0500",x"0800",x"0000",x"FCFF",x"0000",x"FFFF",x"0300",x"0400",x"0200",x"0300",x"FFFF",x"FFFF",x"FBFF",x"F3FF",x"F8FF",x"FCFF",x"0100",x"0600",x"0500",x"0000",x"FDFF",x"FBFF",x"F9FF",x"F9FF",x"FBFF",x"FEFF",x"FEFF",x"0200",x"0200",x"0000",x"0200",x"0100",x"0300",x"0200",x"0300",x"0100",x"0400",x"0300",x"0000",x"FEFF",x"FEFF",x"FDFF",x"FCFF",x"FBFF",x"F4FF",x"F4FF",x"F5FF",x"FCFF",x"FCFF",x"FAFF",x"FDFF",x"FFFF",x"FFFF",x"0200",x"0000",x"0100",x"0300",x"0200",x"0500",x"0500",x"0800",x"0700",x"0600",x"0600",x"0400",x"0400",x"0200",x"0300",x"0300",x"0200",x"0400",x"0400",x"0500",x"0500",x"0300",x"FDFF",x"FEFF",x"0200",x"FFFF",x"0000",x"FDFF",x"FCFF",x"FFFF",x"0100",x"0000",x"0200",x"0500",x"0400",x"0100",x"FEFF",x"FFFF",x"FCFF",x"FEFF",x"0100",x"0000",x"FFFF",x"FEFF",x"FCFF",x"FDFF",x"FBFF",x"FCFF",x"FDFF",x"FEFF",x"0400",x"0700",x"0300",x"0100",x"FEFF",x"FAFF",x"FAFF",x"FBFF",x"FBFF",x"0000",x"0500",x"0200",x"FFFF",x"FBFF",x"FBFF",x"FAFF",x"FEFF",x"0000",x"FCFF",x"FBFF",x"FAFF",x"FBFF",x"FDFF",x"FCFF",x"FDFF",x"0100",x"0100",x"0300",x"0200",x"FFFF",x"FCFF",x"0100",x"0300",x"0600",x"0700",x"0500",x"0800",x"0A00",x"0A00",x"0800",x"0800",x"0A00",x"0A00",x"0100",x"F7FF",x"F6FF",x"F8FF",x"F4FF",x"F4FF",x"FBFF",x"FBFF",x"FAFF",x"FDFF",x"0500",x"0800",x"0900",x"0B00",x"0B00",x"0800",x"0400",x"0000",x"FDFF",x"FCFF",x"FBFF",x"FCFF",x"FFFF",x"0000",x"0300",x"0500",x"0000",x"0400",x"FEFF",x"FEFF",x"0400",x"0200",x"FEFF",x"FEFF",x"0000",x"FBFF",x"FBFF",x"0100",x"0200",x"0100",x"0000",x"FFFF",x"FCFF",x"FEFF",x"FEFF",x"FDFF",x"0100",x"0300",x"0400",x"0800",x"0700",x"0700",x"0600",x"FFFF",x"FFFF",x"0200",x"0200",x"FFFF",x"FDFF",x"FCFF",x"FDFF",x"0100",x"0400",x"0600",x"0700",x"0700",x"0700",x"0700",x"0700",x"0300",x"FDFF",x"FDFF",x"FAFF",x"F6FF",x"F3FF",x"F2FF",x"F2FF",x"F4FF",x"F7FF",x"F6FF",x"F6FF",x"F3FF",x"F3FF",x"F4FF",x"FAFF",x"0000",x"0500",x"0800",x"0900",x"0C00",x"0800",x"0800",x"0E00",x"0E00",x"0D00",x"0C00",x"0700",x"0200",x"FCFF",x"F3FF",x"F3FF",x"EFFF",x"ECFF",x"EAFF",x"EEFF",x"EFFF",x"EFFF",x"F4FF",x"FAFF",x"0D00",x"1500",x"1200",x"1800",x"1D00",x"1B00",x"1900",x"1400",x"1600",x"1300",x"1500",x"0D00",x"0D00",x"0F00",x"0400",x"FEFF",x"F4FF",x"F0FF",x"EAFF",x"E0FF",x"DEFF",x"E0FF",x"E0FF",x"DFFF",x"E2FF",x"EAFF",x"F3FF",x"F6FF",x"FBFF",x"0000",x"0500",x"0800",x"0F00",x"1B00",x"2200",x"2800",x"2B00",x"3100",x"2900",x"1D00",x"1200",x"0900",x"FCFF",x"EBFF",x"E4FF",x"D7FF",x"C8FF",x"BBFF",x"BEFF",x"C2FF",x"C7FF",x"CDFF",x"D5FF",x"E1FF",x"E1FF",x"E6FF",x"F3FF",x"FEFF",x"0A00",x"1200",x"2A00",x"3400",x"4100",x"5000",x"6800",x"8500",x"8F00",x"8E00",x"7C00",x"5D00",x"2C00",x"F1FF",x"B9FF",x"95FF",x"83FF",x"7AFF",x"77FF",x"8DFF",x"A0FF",x"A6FF",x"BBFF",x"CDFF",x"CEFF",x"C1FF",x"BEFF",x"BCFF",x"C0FF",x"E1FF",x"1300",x"6400",x"BF00",x"0E01",x"4F01",x"7D01",x"8901",x"6A01",x"1E01",x"A600",x"1500",x"81FF",x"04FF",x"9FFE",x"5EFE",x"3DFE",x"59FE",x"91FE",x"BAFE",x"DFFE",x"09FF",x"34FF",x"50FF",x"53FF",x"3EFF",x"16FF",x"EFFE",x"E9FE",x"49FF",x"3C00",x"BB01",x"8303",x"3705",x"5206",x"5906",x"3805",x"2503",x"9200",x"08FE",x"04FC",x"D7FA",x"8BFA",x"EDFA",x"A8FB",x"A1FC",x"A0FD",x"74FE",x"3DFF",x"BFFF",x"0B00",x"2700",x"C2FF",x"FAFE",x"FCFD",x"37FD",x"39FD",x"B5FE",x"B001",x"4305",x"7C08",x"9E0A",x"E60A",x"0609",x"D105",x"3F02",x"2CFF",x"D3FC",x"6DFB",x"0BFB",x"58FB",x"1EFC",x"C4FC",x"56FD",x"E4FD",x"BCFE",x"93FF",x"C8FF",x"9DFF",x"C3FE",x"31FD",x"5EFB",x"FFF9",x"D9F8",x"09F8",x"72F8",x"90FA",x"B2FF",x"E106",x"5E0D",x"7F11",x"9712",x"3A10",x"780A",x"8A03",x"97FD",x"B9F9",x"1DF8",x"07F8",x"46F9",x"8DFC",x"AC00",x"4303",x"4D04",x"6304",x"9B03",x"9201",x"61FF",x"0EFD",x"FCF9",x"D8F6",x"7DF4",x"07F4",x"23F5",x"00F7",x"A2F8",x"96F9",x"3FFA",x"3CFA",x"55FD",x"A705",x"C00E",x"0815",x"7E17",x"7516",x"E210",x"8F07",x"59FE",x"0CF8",x"83F5",x"94F5",x"4DF7",x"80FA",x"23FE",x"8A01",x"4604",x"4206",x"3707",x"7A06",x"C404",x"F001",x"F4FD",x"EEF9",x"66F6",x"74F4",x"12F4",x"66F4",x"6CF5",x"73F6",x"47F7",x"A2F7",x"7AF8",x"DDF8",x"02FA",x"5302",x"D40E",x"FB18",x"D81D",x"BA1D",x"C218",x"2E0E",x"F401",x"1BF9",x"37F5",x"DBF4",x"B9F5",x"3DF8",x"C4FB",x"39FF",x"7C02",x"6F04",x"7E05",x"E205",x"B904",x"CE02",x"0A00",x"62FB",x"50F6",x"90F2",x"B9F0",x"61F0",x"6CF1",x"3FF3",x"4EF5",x"9AF6",x"33F7",x"B8F6",x"00F8",x"7502",x"FC11",x"501E",x"6224",x"9124",x"9B1E",x"B811",x"FD01",x"4BF6",x"28F1",x"25F1",x"19F3",x"5DF6",x"71FA",x"A6FD",x"7A00",x"2403",x"FE04",x"9206",x"3707",x"1A06",x"7D02",x"51FC",x"37F6",x"91F0",x"97ED",x"80ED",x"E1EE",x"73F1",x"7AF4",x"94F5",x"01F6",x"79F5",x"4CF4",x"B4FD",x"E510",x"7822",x"3A2C",x"1D2E",x"4428",x"BA19",x"A005",x"55F5",x"5CED",x"98EC",x"5AEF",x"CDF3",x"BCF8",x"76FC",x"D3FE",x"2301",x"3B05",x"CE07",x"7308",x"7D08",x"BD05",x"BFFE",x"97F5",x"E6EE",x"8BEB",x"37EB",x"C9ED",x"9AF0",x"EEF2",x"C0F4",x"5FF4",x"F3F3",x"9EF3",x"C0F8",x"620B",x"AB21",x"E82F",x"E833",x"222F",x"A521",x"550C",x"81F7",x"63EB",x"00E8",x"49EB",x"BBF0",x"A2F6",x"0CFC",x"57FF",x"AB01",x"3B06",x"D109",x"B809",x"A707",x"FB04",x"5EFF",x"B0F6",x"1BF0",x"18EB",x"34EA",x"B4EA",x"A7EE",x"B1F1",x"88F2",x"ACF3",x"A9F3",x"41F3",x"7DF5",x"7F05",x"3C1D",x"5C2F",x"FC35",x"2233",x"1B28",x"F213",x"6AFC",x"D9EC",x"03E7",x"A3E8",x"DCED",x"34F4",x"B9FB",x"5F01",x"5903",x"1304",x"4005",x"4605",x"A903",x"6D02",x"9B01",x"7EFD",x"73F5",x"22EF",x"46ED",x"17EB",x"61EC",x"7EEE",x"A9F1",x"E5F2",x"58F4",x"42F5",x"14F6",x"4B04",x"BE1C",x"B530",x"1139",x"4536",x"5B2A",x"2915",x"99FC",x"32EA",x"49E2",x"FCE4",x"18EC",x"95F4",x"8BFC",x"3102",x"0A05",x"6F04",x"4704",x"C804",x"3405",x"9E04",x"A101",x"53FB",x"B0F3",x"8CEE",x"02EB",x"1AEB",x"D7ED",x"5FF0",x"28F2",x"95F2",x"85F1",x"80F2",x"59F2",x"BF00",x"E91E",x"1038",x"D03F",x"8238",x"DE28",x"6111",x"DAF6",x"17E4",x"29DF",x"DFE5",x"28F1",x"A0FA",x"D001",x"B203",x"7A01",x"BB01",x"C703",x"2D04",x"5104",x"5405",x"A701",x"49FA",x"1DF1",x"C8EA",x"AEE9",x"93EC",x"DEEE",x"D9EF",x"13F2",x"50F1",x"D9F0",x"05F1",x"60F2",x"3108",x"472C",x"7644",x"0545",x"9234",x"691D",x"CF03",x"95EB",x"29DE",x"D8E0",x"57EE",x"D8FA",x"F200",x"8502",x"EAFF",x"28FB",x"5FFC",x"E603",x"A609",x"0F0B",x"3009",x"DD02",x"AAF7",x"82EC",x"76E6",x"2EE6",x"8FEA",x"62F0",x"6BF3",x"E8F1",x"EBEB",x"70E9",x"3EE7",x"C8F0",x"EA17",x"6744",x"4656",x"8B46",x"B927",x"9E09",x"83F1",x"35E2",x"17E2",x"31F1",x"0F03",x"530A",x"A805",x"9CFB",x"E8F1",x"C9ED",x"45F8",x"AB0A",x"DC14",x"0E13",x"AB09",x"EBFB",x"D6EA",x"D6DE",x"7EDE",x"FFE6",x"34F1",x"B6F6",x"C6F4",x"A9ED",x"E0E4",x"53E0",x"62E0",x"4BFE",x"3B3A",x"3F65",x"4D5D",x"B530",x"0905",x"78EB",x"A4E1",x"48E4",x"07F5",x"E10B",x"FA15",x"6A0A",x"2BF6",x"D2E7",x"8AE4",x"95F1",x"A40D",x"F821",x"371F",x"CE0D",x"FEFA",x"08EA",x"ACDD",x"A5DD",x"E4E8",x"4AF4",x"B5F8",x"A0F3",x"5FEA",x"6FE0",x"08DC",x"16DC",x"61F2",x"0B31",x"D368",x"1966",x"2F31",x"B0FE",x"04E9",x"E8E8",x"8CF0",x"67FF",x"9111",x"2F16",x"2703",x"E8E9",x"72DF",x"86E6",x"1CF6",x"010C",x"4322",x"1A22",x"0A0C",x"F7F7",x"0CEF",x"4DE9",x"30E6",x"F6EB",x"FCF3",x"C9F4",x"0AEF",x"E2E7",x"DFE0",x"E6DC",x"D1DD",x"3AE7",x"E11A",x"985C",x"5368",x"C635",x"B5FE",x"B4EC",x"BEF4",x"A5FC",x"B403",x"4B10",x"F813",x"F500",x"C1E6",x"5DDF",x"4CEA",x"B3F9",x"1C07",x"A814",x"C61B",x"F310",x"D1FD",x"4BF4",x"29F1",x"2CEC",x"4CEB",x"E8F0",x"A1F4",x"1BF1",x"5EE8",x"AFE2",x"93DE",x"6BE1",x"A6E2",x"39FB",x"113D",x"0A66",x"FC48",x"E10C",x"33F2",x"82FB",x"5F05",x"2704",x"F109",x"1613",x"6009",x"E4EE",x"96E2",x"C2EC",x"A1F9",x"9BFE",x"0903",x"6511",x"3319",x"370C",x"27FB",x"6FF3",x"6CEF",x"F9EA",x"76ED",x"74F3",x"20F3",x"58ED",x"04E8",x"0FE4",x"D7DF",x"6AE1",x"6AE6",x"8412",x"2A54",x"455F",x"832B",x"2CFC",x"ECF8",x"0B05",x"9602",x"B200",x"D00C",x"0510",x"8FFB",x"E9E5",x"A6E8",x"3DF6",x"23FB",x"F1FD",x"F308",x"7213",x"BE10",x"6006",x"1EFD",x"C6F4",x"12ED",x"DDEB",x"1FF2",x"13F7",x"7DF4",x"80EB",x"99E2",x"92DD",x"BBDE",x"18E5",x"70ED",x"8D1F",x"015A",x"D253",x"171B",x"87F9",x"DD01",x"CD0A",x"D103",x"7205",x"4F11",x"580A",x"7DEF",x"98E1",x"E6EC",x"D1F7",x"61F9",x"2DFF",x"C70A",x"E312",x"F812",x"9809",x"00FB",x"37F0",x"F7EF",x"12F6",x"54F9",x"CCF7",x"E7F0",x"99E6",x"D1DC",x"1BD9",x"A6DE",x"03EC",x"0BF9",x"F21C",x"F946",x"C345",x"3D20",x"4606",x"5208",x"520B",x"9B05",x"E406",x"7D0C",x"4301",x"FEEB",x"65E5",x"FAF0",x"F1FA",x"3EFD",x"3300",x"4E04",x"E807",x"BB0E",x"5112",x"2A06",x"C4F4",x"1FF2",x"25F9",x"4AF9",x"92F2",x"3CEB",x"75E4",x"E8DD",x"42DE",x"0DE5",x"74F0",x"FBEB",x"70F5",x"703F",x"C86A",x"7C3A",x"3300",x"B400",x"030F",x"0401",x"41F9",x"D209",x"0408",x"9EEA",x"8BDD",x"A7F0",x"6A00",x"48FC",x"90FB",x"4D02",x"F602",x"8D06",x"4514",x"3416",x"4703",x"79F2",x"4FF3",x"C9F9",x"4AF9",x"82F2",x"3AE8",x"34E0",x"71E0",x"F9E6",x"C5ED",x"E7F3",x"A7ED",x"3EFA",x"6B41",x"E961",x"1F32",x"DE06",x"9E0A",x"0708",x"CBF3",x"02FA",x"410D",x"1600",x"EEE6",x"B6E6",x"FAF5",x"85FC",x"42FB",x"0AFF",x"3700",x"C901",x"A809",x"1218",x"9C19",x"5904",x"F4F2",x"F5F1",x"A5F6",x"B2F4",x"00EE",x"9BE8",x"CFE4",x"ABE3",x"2AE8",x"8DF0",x"F7F7",x"69EF",x"57EE",x"0635",x"BA61",x"FA36",x"EC0F",x"9D0E",x"0FFD",x"19E7",x"97FB",x"D913",x"0701",x"77E8",x"FFE8",x"A1EE",x"4EF6",x"FE00",x"0C06",x"2303",x"3706",x"290F",x"8F10",x"E30F",x"E50A",x"0AF9",x"48ED",x"A0EF",x"62F1",x"C5EF",x"13ED",x"51E8",x"05E6",x"88E8",x"D1F1",x"CFF8",x"19F5",x"8AEF",x"C325",x"BE55",x"DE39",x"AA19",x"0A0E",x"78F7",x"39EA",x"5201",x"680E",x"3FFC",x"C3EC",x"68EB",x"C4EA",x"AFF5",x"C203",x"5A07",x"3706",x"5107",x"8A07",x"FD12",x"9D18",x"DA0B",x"73F9",x"BBEC",x"E7EC",x"61F2",x"8DF4",x"5CEF",x"03E7",x"0CE6",x"05E9",x"F3F1",x"EAFB",x"D7FB",x"3FEF",x"580C",x"E145",x"AD3C",x"D11F",x"8315",x"D600",x"1EED",x"16F9",x"EB05",x"07FF",x"2FF5",x"0AEF",x"FEE6",x"34F1",x"5203",x"B408",x"0108",x"3D0A",x"1D0E",x"1C0E",x"4A10",x"D80B",x"D9FB",x"C3EE",x"14ED",x"E0EF",x"DEF2",x"81F1",x"92EB",x"0DE9",x"10EC",x"63F0",x"8CFB",x"6201",x"CEFA",x"25F2",x"F417",x"9B3B",x"8C2D",x"3923",x"2816",x"B6F8",x"80F0",x"39FE",x"EDFF",x"2CFB",x"E8F7",x"F2EE",x"FFEB",x"35FB",x"BB03",x"EF04",x"160A",x"650D",x"A80D",x"540F",x"140D",x"D202",x"88F5",x"FAED",x"95EF",x"86F2",x"84F2",x"1DEF",x"A6EA",x"7AE9",x"E9EE",x"4FFA",x"A903",x"6002",x"CCFD",x"9BFC",x"E60F",x"8F21",x"1025",x"DE23",x"1C15",x"1D03",x"3BFD",x"FDFB",x"FAF7",x"89F6",x"4CF5",x"F0F3",x"99F7",x"2CFD",x"7BFE",x"E200",x"7804",x"1508",x"1E0B",x"0B0E",x"440C",x"2303",x"D1F9",x"A1F3",x"D7F0",x"96F1",x"F4F3",x"71F5",x"CCF3",x"A4F2",x"33F6",x"B8FA",x"77FD",x"32FF",x"8CFF",x"F6FD",x"A6FC",x"E907",x"D310",x"5113",x"3E17",x"6317",x"3314",x"E60D",x"F805",x"54FC",x"D4F3",x"75F0",x"E8F0",x"56F3",x"02FA",x"E1FF",x"3B03",x"8504",x"2F07",x"1F09",x"EC07",x"EC06",x"4504",x"8AFE",x"29F9",x"50F4",x"A8F0",x"0FF1",x"E2F2",x"26F4",x"1EF7",x"17FB",x"90FD",x"90FD",x"1AFD",x"94FD",x"A2FD",x"D800",x"1409",x"2A0E",x"5D12",x"1B16",x"F813",x"0910",x"AD0C",x"6305",x"B2FC",x"A8F6",x"57F3",x"60F4",x"E1F6",x"DCF8",x"7AFB",x"CFFF",x"9902",x"1803",x"E205",x"BF07",x"1606",x"2003",x"87FF",x"65FA",x"ACF6",x"A5F4",x"CAF3",x"7AF4",x"76F7",x"82FA",x"0AFB",x"ACFA",x"8FFB",x"DAFB",x"94FB",x"09FE",x"9B03",x"5A09",x"D50D",x"F513",x"0317",x"4815",x"5010",x"D107",x"ACFF",x"4FFB",x"1FF8",x"DDF5",x"77F5",x"F7F6",x"32FA",x"A9FD",x"8300",x"B303",x"F804",x"6804",x"9904",x"DB04",x"9E02",x"92FD",x"E7F8",x"3EF6",x"E4F4",x"7FF5",x"5BF6",x"2EF7",x"00F8",x"A5F9",x"4CFB",x"2AFC",x"84FD",x"D7FF",x"3702",x"B205",x"DE0B",x"1210",x"9512",x"7C12",x"290E",x"E908",x"8A05",x"F000",x"C4FA",x"7DF7",x"45F7",x"39F7",x"E2F8",x"89FC",x"4B00",x"2702",x"0902",x"DA02",x"BB03",x"5A04",x"A102",x"69FF",x"62FC",x"D6F8",x"64F6",x"63F6",x"E3F5",x"30F6",x"FDF8",x"06FA",x"4FFB",x"93FD",x"A4FE",x"5AFF",x"BB00",x"0003",x"5206",x"2409",x"AD0C",x"F90D",x"8F0D",x"4B0C",x"C008",x"0F05",x"5601",x"E0FE",x"B9FC",x"D2F9",x"7EFA",x"CFFC",x"9BFD",x"41FF",x"8400",x"8001",x"0802",x"4402",x"5101",x"5EFF",x"C6FC",x"47FA",x"83F9",x"2AF9",x"55F8",x"BEF7",x"EBF8",x"35FA",x"8CFB",x"44FE",x"3EFF",x"4DFF",x"5000",x"0A01",x"B502",x"5505",x"DC07",x"D109",x"570A",x"190A",x"8E08",x"6806",x"6604",x"B401",x"D9FE",x"B5FD",x"B9FD",x"99FD",x"5DFD",x"9EFD",x"61FE",x"C3FE",x"B9FF",x"3800",x"48FF",x"3CFE",x"B3FC",x"7CFB",x"71FB",x"CCFA",x"57FA",x"27FA",x"66FA",x"C0FB",x"25FD",x"C9FD",x"EAFD",x"CCFE",x"0000",x"2A01",x"DA01",x"D303",x"8904",x"5C05",x"E206",x"5007",x"5907",x"FD06",x"FD04",x"6C03",x"1E02",x"4C01",x"6100",x"89FF",x"FDFE",x"3DFE",x"06FF",x"36FF",x"A4FF",x"6CFF",x"1CFE",x"6EFD",x"84FD",x"18FD",x"C4FC",x"7AFC",x"15FC",x"74FB",x"BDFB",x"9CFC",x"02FD",x"59FD",x"C7FE",x"2BFF",x"D0FF",x"7B00",x"0901",x"E401",x"1E02",x"9702",x"0303",x"E603",x"0004",x"F703",x"AA03",x"F402",x"9C03",x"DF02",x"9201",x"A900",x"BBFF",x"93FF",x"8000",x"0201",x"9700",x"CAFF",x"31FF",x"28FF",x"9DFF",x"97FF",x"B9FE",x"14FE",x"3DFD",x"02FD",x"CEFC",x"46FC",x"E3FB",x"7BFC",x"D5FC",x"6EFD",x"C3FE",x"B6FF",x"4A00",x"9C00",x"A300",x"F400",x"A101",x"E301",x"D801",x"3C01",x"C300",x"7101",x"8F01",x"6402",x"1202",x"BE01",x"8401",x"6601",x"DF01",x"9701",x"C600",x"5500",x"0900",x"0D00",x"5E00",x"1600",x"F7FF",x"5EFF",x"24FF",x"C2FE",x"7FFE",x"0BFE",x"46FE",x"00FE",x"90FD",x"28FE",x"99FE",x"B0FE",x"9FFE",x"AEFE",x"48FF",x"E9FF",x"C700",x"EF00",x"E000",x"EA00",x"DA00",x"1501",x"8501",x"7101",x"5D01",x"C400",x"6200",x"D200",x"4101",x"F500",x"DC00",x"B500",x"C300",x"0B01",x"D300",x"D900",x"9900",x"4600",x"1300",x"ACFF",x"75FF",x"8BFF",x"B4FE",x"62FE",x"84FE",x"1FFE",x"0BFE",x"41FE",x"9AFE",x"DDFE",x"00FF",x"8DFF",x"E0FF",x"ECFF",x"D2FF",x"A6FF",x"0000",x"9300",x"8600",x"A500",x"5700",x"1700",x"A800",x"0301",x"4101",x"1D01",x"B300",x"4E00",x"1700",x"1300",x"3E00",x"7E00",x"9E00",x"E300",x"D800",x"7A00",x"3200",x"ADFF",x"4BFF",x"2CFF",x"2FFF",x"0AFF",x"FFFE",x"11FF",x"B0FE",x"E9FE",x"BBFF",x"0300",x"1200",x"FAFF",x"0700",x"2F00",x"3500",x"4A00",x"4C00",x"6700",x"4900",x"3600",x"8300",x"C300",x"8000",x"7000",x"6700",x"5800",x"6200",x"4400",x"4700",x"4800",x"3000",x"6B00",x"5700",x"0C00",x"ACFF",x"5CFF",x"73FF",x"A5FF",x"AEFF",x"8AFF",x"5BFF",x"37FF",x"13FF",x"53FF",x"B6FF",x"F6FF",x"2900",x"2800",x"2200",x"2600",x"4700",x"1400",x"1900",x"4C00",x"5100",x"6B00",x"5500",x"1200",x"E3FF",x"D5FF",x"EEFF",x"2300",x"2A00",x"5000",x"7700",x"8F00",x"9000",x"6700",x"1400",x"C5FF",x"84FF",x"5EFF",x"90FF",x"7AFF",x"3EFF",x"42FF",x"33FF",x"60FF",x"B9FF",x"FDFF",x"3900",x"4100",x"1500",x"0A00",x"0100",x"1300",x"0F00",x"3C00",x"6C00",x"5700",x"3200",x"1400",x"FDFF",x"0000",x"2C00",x"5E00",x"8800",x"9500",x"6000",x"3900",x"4200",x"4A00",x"4A00",x"4B00",x"3000",x"F9FF",x"D2FF",x"B3FF",x"B1FF",x"A8FF",x"8DFF",x"ABFF",x"9CFF",x"AFFF",x"E9FF",x"F1FF",x"FDFF",x"0A00",x"1A00",x"3B00",x"4000",x"4300",x"4500",x"2A00",x"0600",x"F2FF",x"E3FF",x"C1FF",x"B6FF",x"D1FF",x"FBFF",x"FEFF",x"1B00",x"2700",x"2B00",x"3700",x"1D00",x"1800",x"2200",x"0A00",x"F0FF",x"D5FF",x"B8FF",x"ABFF",x"A0FF",x"98FF",x"ABFF",x"B3FF",x"B6FF",x"EEFF",x"1100",x"1D00",x"1900",x"2800",x"3600",x"3400",x"2000",x"0900",x"F0FF",x"F4FF",x"FCFF",x"FCFF",x"0400",x"1000",x"0800",x"FFFF",x"FDFF",x"0100",x"1800",x"2D00",x"3000",x"3800",x"3400",x"2D00",x"3500",x"2700",x"0F00",x"FBFF",x"F6FF",x"F1FF",x"EBFF",x"E1FF",x"D5FF",x"D3FF",x"E7FF",x"EBFF",x"ECFF",x"FBFF",x"FFFF",x"0100",x"FCFF",x"F2FF",x"F4FF",x"E6FF",x"D5FF",x"E3FF",x"0100",x"1500",x"0B00",x"0300",x"0200",x"0000",x"2400",x"4500",x"3E00",x"3100",x"1400",x"FDFF",x"FDFF",x"0500",x"1900",x"1A00",x"FFFF",x"FFFF",x"FAFF",x"FAFF",x"0C00",x"FFFF",x"E9FF",x"E2FF",x"EBFF",x"F2FF",x"F5FF",x"F3FF",x"D7FF",x"C6FF",x"CAFF",x"DEFF",x"F5FF",x"0000",x"FDFF",x"FFFF",x"0200",x"1000",x"0F00",x"0C00",x"0A00",x"0C00",x"1C00",x"2500",x"1F00",x"1400",x"FFFF",x"ECFF",x"F0FF",x"0900",x"0E00",x"0600",x"0600",x"FDFF",x"FFFF",x"0200",x"0000",x"F6FF",x"EDFF",x"E9FF",x"F2FF",x"F9FF",x"0300",x"FBFF",x"E7FF",x"DCFF",x"E6FF",x"F9FF",x"FBFF",x"F6FF",x"F0FF",x"E1FF",x"E5FF",x"FCFF",x"0D00",x"1300",x"1C00",x"1C00",x"2400",x"2E00",x"2900",x"1700",x"0900",x"0700",x"1700",x"2300",x"2200",x"1E00",x"0800",x"FEFF",x"FDFF",x"0800",x"1200",x"0000",x"E8FF",x"DEFF",x"D9FF",x"EAFF",x"F2FF",x"F2FF",x"F2FF",x"F6FF",x"FBFF",x"F7FF",x"F6FF",x"F9FF",x"F5FF",x"0400",x"1200",x"1000",x"EEFF",x"ECFF",x"EFFF",x"1500",x"CB00",x"A100",x"4400",x"DAFF",x"5AFF",x"58FF",x"89FF",x"CBFF",x"1900",x"3100",x"3100",x"0000",x"E2FF",x"D1FF",x"BCFF",x"D4FF",x"E2FF",x"FEFF",x"1600",x"0C00",x"0E00",x"FCFF",x"FAFF",x"1200",x"2D00",x"3300",x"0E00",x"F3FF",x"EEFF",x"E1FF",x"FDFF",x"2900",x"3900",x"3D00",x"2100",x"0200",x"E9FF",x"E6FF",x"0800",x"1C00",x"2100",x"2900",x"2200",x"0900",x"EDFF",x"EDFF",x"F8FF",x"0400",x"2000",x"1F00",x"0800",x"ECFF",x"DEFF",x"DBFF",x"EDFF",x"0F00",x"2300",x"2100",x"1900",x"FFFF",x"F4FF",x"E3FF",x"E2FF",x"F1FF",x"F6FF",x"0E00",x"1500",x"0D00",x"0100",x"EBFF",x"DCFF",x"EAFF",x"FBFF",x"0100",x"0400",x"0500",x"F5FF",x"F1FF",x"E8FF",x"EAFF",x"FAFF",x"FBFF",x"FAFF",x"F7FF",x"FCFF",x"F9FF",x"F2FF",x"EDFF",x"ECFF",x"E9FF",x"F0FF",x"0F00",x"1000",x"0A00",x"1800",x"1200",x"0900",x"0F00",x"F8FF",x"E5FF",x"F1FF",x"F2FF",x"FBFF",x"1000",x"0400",x"EDFF",x"FBFF",x"0500",x"F7FF",x"0F00",x"2700",x"0900",x"0500",x"1900",x"0A00",x"FCFF",x"0A00",x"FAFF",x"E5FF",x"0100",x"1300",x"0E00",x"0300",x"FAFF",x"F1FF",x"F3FF",x"0700",x"1900",x"0300",x"FCFF",x"0600",x"1100",x"0E00",x"0A00",x"1200",x"0400",x"0200",x"0200",x"F8FF",x"EFFF",x"E8FF",x"F1FF",x"FAFF",x"F9FF",x"0C00",x"0F00",x"0900",x"0700",x"0800",x"FDFF",x"FAFF",x"0D00",x"0E00",x"FFFF",x"FCFF",x"F7FF",x"EFFF",x"FBFF",x"0900",x"0D00",x"0500",x"F7FF",x"F0FF",x"F0FF",x"F0FF",x"FFFF",x"1100",x"2000",x"2300",x"0600",x"EDFF",x"E1FF",x"E0FF",x"E5FF",x"F0FF",x"F9FF",x"F6FF",x"FEFF",x"0200",x"FCFF",x"0600",x"1200",x"1200",x"1000",x"0900",x"0300",x"FDFF",x"F6FF",x"F4FF",x"F9FF",x"0300",x"0D00",x"0D00",x"0D00",x"0200",x"F2FF",x"F5FF",x"FBFF",x"FBFF",x"FBFF",x"0200",x"0300",x"0100",x"FDFF",x"F9FF",x"F5FF",x"F9FF",x"FBFF",x"FDFF",x"FCFF",x"EEFF",x"EFFF",x"FCFF",x"0200",x"0C00",x"1000",x"0900",x"0800",x"0F00",x"0E00",x"0A00",x"1300",x"1200",x"0500",x"FFFF",x"FCFF",x"FAFF",x"0200",x"0800",x"0500",x"0500",x"0500",x"F8FF",x"FCFF",x"0200",x"0600",x"0B00",x"0900",x"0C00",x"0A00",x"0200",x"F8FF",x"EDFF",x"F3FF",x"F4FF",x"F2FF",x"F9FF",x"FBFF",x"FCFF",x"FFFF",x"FBFF",x"F8FF",x"FBFF",x"0300",x"0900",x"0C00",x"0D00",x"0900",x"FFFF",x"F9FF",x"F6FF",x"F4FF",x"F6FF",x"FAFF",x"0100",x"FDFF",x"F6FF",x"F6FF",x"F7FF",x"F7FF",x"FBFF",x"0500",x"0700",x"0300",x"0100",x"0200",x"0100",x"0200",x"0100",x"0500",x"0700",x"0600",x"0500",x"FEFF",x"FCFF",x"F9FF",x"FDFF",x"0100",x"0000",x"FCFF",x"F7FF",x"F7FF",x"F6FF",x"F9FF",x"0200",x"0200",x"0400",x"FEFF",x"F8FF",x"FEFF",x"0500",x"0A00",x"0D00",x"0D00",x"0A00",x"0700",x"0800",x"0800",x"0C00",x"0D00",x"0D00",x"0A00",x"0400",x"FEFF",x"FAFF",x"F9FF",x"F4FF",x"F5FF",x"F4FF",x"F7FF",x"FAFF",x"FFFF",x"0100",x"0300",x"0200",x"0300",x"0700",x"0400",x"0300",x"0800",x"0B00",x"0600",x"0700",x"0700",x"0600",x"0400",x"0600",x"0300",x"0100",x"0200",x"F8FF",x"F3FF",x"F3FF",x"F3FF",x"F6FF",x"F6FF",x"F8FF",x"FCFF",x"FEFF",x"FFFF",x"FEFF",x"FDFF",x"F9FF",x"FAFF",x"FDFF",x"0200",x"0200",x"0100",x"0200",x"0200",x"F9FF",x"F8FF",x"FBFF",x"FEFF",x"FDFF",x"FEFF",x"FEFF",x"FEFF",x"FDFF",x"FBFF",x"FCFF",x"F8FF",x"FEFF",x"FCFF",x"FAFF",x"FEFF",x"FAFF",x"FDFF",x"0200",x"0700",x"0700",x"0700",x"0900",x"0800",x"0800",x"0B00",x"0800",x"0800",x"0700",x"0200",x"FDFF",x"F9FF",x"FAFF",x"FAFF",x"FDFF",x"0100",x"0200",x"FCFF",x"FDFF",x"F9FF",x"FBFF",x"0400",x"0B00",x"1000",x"1000",x"0F00",x"0C00",x"0B00",x"0B00",x"0B00",x"0F00",x"1200",x"0C00",x"0700",x"0200",x"F9FF",x"F9FF",x"FAFF",x"FBFF",x"FFFF",x"FEFF",x"FDFF",x"FBFF",x"F5FF",x"F1FF",x"F0FF",x"F0FF",x"F2FF",x"F7FF",x"F8FF",x"F7FF",x"F7FF",x"F6FF",x"F5FF",x"F5FF",x"F9FF",x"FBFF",x"FCFF",x"FBFF",x"F9FF",x"FBFF",x"0000",x"0500",x"0900",x"0800",x"0700",x"0400",x"FEFF",x"FDFF",x"FAFF",x"FCFF",x"FEFF",x"FEFF",x"FEFF",x"F9FF",x"F8FF",x"FAFF",x"FFFF",x"0400",x"0700",x"0700",x"0C00",x"0D00",x"0B00",x"0900",x"0700",x"0700",x"0B00",x"0A00",x"0800",x"0400",x"0200",x"0100",x"FCFF",x"F9FF",x"F9FF",x"FBFF",x"FDFF",x"FDFF",x"0100",x"0500",x"0900",x"0B00",x"0D00",x"0C00",x"0800",x"0900",x"0500",x"0500",x"0900",x"0600",x"0300",x"0200",x"0300",x"0200",x"0100",x"0300",x"0100",x"0100",x"0100",x"0100",x"FFFF",x"FBFF",x"FAFF",x"FAFF",x"FAFF",x"FAFF",x"FAFF",x"F8FF",x"F7FF",x"FAFF",x"F9FF",x"FAFF",x"FEFF",x"FDFF",x"FAFF",x"FAFF",x"FAFF",x"FDFF",x"FDFF",x"F9FF",x"F7FF",x"F5FF",x"F5FF",x"F7FF",x"F6FF",x"F8FF",x"F9FF",x"FAFF",x"FCFF",x"FFFF",x"0100",x"0100",x"0100",x"0100",x"0100",x"0100",x"0100",x"0200",x"FFFF",x"0000",x"0200",x"0200",x"0000",x"0000",x"0100",x"0200",x"0500",x"0800",x"0700",x"0900",x"0A00",x"0500",x"0300",x"0400",x"0500",x"0700",x"0900",x"0700",x"0500",x"0600",x"0700",x"0900",x"0800",x"0A00",x"0A00",x"0A00",x"0A00",x"0400",x"0100",x"0000",x"FFFF",x"FEFF",x"FEFF",x"FCFF",x"F8FF",x"F6FF",x"F5FF",x"F6FF",x"F4FF",x"F7FF",x"FBFF",x"FAFF",x"F7FF",x"F7FF",x"F8FF",x"FBFF",x"FFFF",x"0200",x"0800",x"0B00",x"0800",x"0600",x"0300",x"0300",x"0100",x"FFFF",x"FEFF",x"0200",x"0200",x"0100",x"0000",x"0000",x"0200",x"F8FF",x"F8FF",x"FAFF",x"F9FF",x"FAFF",x"FAFF",x"F9FF",x"F8FF",x"FCFF",x"FCFF",x"FAFF",x"FEFF",x"FFFF",x"FEFF",x"FFFF",x"FFFF",x"0200",x"0200",x"0200",x"0100",x"0000",x"0000",x"0100",x"0400",x"0200",x"0500",x"0900",x"0700",x"0800",x"0600",x"0500",x"0500",x"0300",x"0100",x"FCFF",x"FAFF",x"FAFF",x"FBFF",x"FFFF",x"0400",x"0700",x"0300",x"FFFF",x"FEFF",x"FBFF",x"FAFF",x"FAFF",x"FCFF",x"FDFF",x"FBFF",x"FAFF",x"FAFF",x"0000",x"0100",x"0400",x"0900",x"0900",x"0C00",x"0E00",x"0C00",x"0800",x"0A00",x"0700",x"0400",x"0600",x"0500",x"0100",x"FEFF",x"FDFF",x"F9FF",x"F6FF",x"F7FF",x"F6FF",x"F8FF",x"FAFF",x"FBFF",x"FCFF",x"FDFF",x"FFFF",x"FFFF",x"0100",x"0000",x"0000",x"0000",x"FEFF",x"FBFF",x"FCFF",x"FCFF",x"FAFF",x"FAFF",x"FBFF",x"FBFF",x"FCFF",x"FCFF",x"FBFF",x"FAFF",x"FAFF",x"FFFF",x"0000",x"FFFF",x"FCFF",x"FFFF",x"FEFF",x"0000",x"0200",x"0200",x"0700",x"0800",x"0600",x"0400",x"0400",x"0200",x"0100",x"0000",x"0300",x"0500",x"0500",x"0300",x"0400",x"0500",x"0600",x"0400",x"0300",x"0100",x"0000",x"FDFF",x"FAFF",x"FBFF",x"FFFF",x"FEFF",x"FFFF",x"0300",x"0200",x"0200",x"FFFF",x"FFFF",x"0400",x"0400",x"0300",x"0200",x"0200",x"FFFF",x"FEFF",x"FFFF",x"0000",x"0300",x"0100",x"0200",x"0300",x"0100",x"0100",x"0200",x"0000",x"0000",x"FDFF",x"FFFF",x"0100",x"0100",x"FEFF",x"FBFF",x"FDFF",x"FDFF",x"FDFF",x"0000",x"0100",x"0000",x"FDFF",x"FDFF",x"FCFF",x"FAFF",x"FFFF",x"0100",x"0100",x"0800",x"0500",x"0500",x"0600",x"0200",x"0200",x"0000",x"0200",x"0200",x"0300",x"0100",x"FEFF",x"FDFF",x"FFFF",x"FCFF",x"FBFF",x"FAFF",x"FAFF",x"FAFF",x"FAFF",x"F8FF",x"F4FF",x"F6FF",x"F9FF",x"F7FF",x"F7FF",x"F9FF",x"FFFF",x"0200",x"0400",x"0300",x"0400",x"0600",x"0400",x"0700",x"0600",x"0700",x"0900",x"0A00",x"0800",x"0500",x"0100",x"0100",x"0100",x"0000",x"0000",x"0100",x"0100",x"0000",x"0100",x"0100",x"0000",x"FFFF",x"0100",x"FFFF",x"0100",x"0300",x"0100",x"FFFF",x"FFFF",x"FEFF",x"FFFF",x"0100",x"0100",x"0300",x"0200",x"0400",x"0400",x"0000",x"0100",x"FEFF",x"FAFF",x"FBFF",x"FCFF",x"FDFF",x"FDFF",x"FDFF",x"FDFF",x"FFFF",x"FCFF",x"FDFF",x"FEFF",x"FFFF",x"FDFF",x"FFFF",x"FFFF",x"FEFF",x"0000",x"0000",x"0000",x"0100",x"0400",x"0000",x"0300",x"0600",x"0600",x"0700",x"0600",x"0700",x"0800",x"0300",x"0200",x"0300",x"0100",x"0000",x"FDFF",x"FEFF",x"FDFF",x"FEFF",x"FCFF",x"FFFF",x"0000",x"0000",x"FEFF",x"FCFF",x"FAFF",x"FDFF",x"FDFF",x"FDFF",x"FCFF",x"FBFF",x"FCFF",x"0000",x"0200",x"FEFF",x"FFFF",x"FFFF",x"FBFF",x"FDFF",x"FEFF",x"0100",x"0200",x"0400",x"0600",x"0400",x"0500",x"0200",x"0300",x"0200",x"0100",x"FFFF",x"0100",x"FCFF",x"F6FF",x"F8FF",x"FAFF",x"F8FF",x"FBFF",x"FFFF",x"FFFF",x"0000",x"FFFF",x"0000",x"0200",x"0200",x"0400",x"0B00",x"0A00",x"0500",x"0400",x"0200",x"0100",x"0100",x"0400",x"0200",x"FFFF",x"FCFF",x"FCFF",x"FEFF",x"FFFF",x"0100",x"0100",x"0400",x"0500",x"0600",x"0700",x"0700",x"0700",x"0500",x"0300",x"0400",x"0200",x"0200",x"0100",x"FEFF",x"0100",x"FDFF",x"FEFF",x"FCFF",x"FAFF",x"FBFF",x"FBFF",x"FAFF",x"FBFF",x"FBFF",x"FAFF",x"F7FF",x"FAFF",x"FCFF",x"FCFF",x"FEFF",x"0200",x"0100",x"0000",x"0000",x"FEFF",x"FAFF",x"F8FF",x"F7FF",x"F8FF",x"FBFF",x"FDFF",x"FAFF",x"FBFF",x"FFFF",x"FCFF",x"FCFF",x"FFFF",x"0000",x"0600",x"0600",x"0500",x"0600",x"0500",x"0500",x"0700",x"0C00",x"0C00",x"0C00",x"1000",x"0B00",x"0700",x"0600",x"0900",x"0A00",x"0900",x"0600",x"0200",x"0300",x"0300",x"0100",x"0000",x"0100",x"FEFF",x"FEFF",x"FCFF",x"FBFF",x"FCFF",x"FAFF",x"F8FF",x"F6FF",x"F8FF",x"F7FF",x"FAFF",x"F9FF",x"F8FF",x"FCFF",x"FDFF",x"F9FF",x"F8FF",x"F6FF",x"F7FF",x"F6FF",x"F7FF",x"F6FF",x"F9FF",x"FDFF",x"FFFF",x"FEFF",x"FEFF",x"FFFF",x"0100",x"0100",x"0200",x"0300",x"0400",x"0600",x"0500",x"0500",x"0500",x"0300",x"0500",x"0700",x"0900",x"0A00",x"0700",x"0800",x"0500",x"0500",x"0300",x"0300",x"0300",x"0100",x"FEFF",x"FEFF",x"FFFF",x"FFFF",x"0400",x"0600",x"0B00",x"0B00",x"0B00",x"0700",x"0300",x"0100",x"FCFF",x"FCFF",x"FDFF",x"FFFF",x"0000",x"FFFF",x"FFFF",x"FEFF",x"0100",x"FCFF",x"FCFF",x"FEFF",x"FEFF",x"FCFF",x"FEFF",x"FFFF",x"FFFF",x"0000",x"0000",x"FEFF",x"FCFF",x"FDFF",x"FFFF",x"0000",x"0300",x"0200",x"FEFF",x"FBFF",x"F8FF",x"FAFF",x"FAFF",x"F8FF",x"F9FF",x"FBFF",x"FEFF",x"FEFF",x"FDFF",x"F9FF",x"FBFF",x"FEFF",x"F9FF",x"F8FF",x"F9FF",x"FCFF",x"FCFF",x"FEFF",x"0200",x"0900",x"0900",x"0700",x"0900",x"0800",x"0300",x"FEFF",x"FFFF",x"FEFF",x"FAFF",x"F9FF",x"FBFF",x"0100",x"FEFF",x"FEFF",x"0000",x"0100",x"0300",x"0400",x"0400",x"0200",x"FEFF",x"FCFF",x"0100",x"0200",x"0300",x"0300",x"0200",x"0500",x"0400",x"0400",x"0300",x"0300",x"0100",x"0100",x"0100",x"0400",x"0300",x"0400",x"0300",x"0300",x"0500",x"0500",x"0700",x"0900",x"0900",x"0700",x"0400",x"0000",x"FCFF",x"FCFF",x"FBFF",x"FEFF",x"FDFF",x"FEFF",x"0000",x"0000",x"0000",x"FFFF",x"FCFF",x"FAFF",x"FEFF",x"FEFF",x"FCFF",x"0000",x"0200",x"0100",x"0000",x"0000",x"FEFF",x"FBFF",x"FDFF",x"FEFF",x"FFFF",x"FCFF",x"FAFF",x"FAFF",x"F9FF",x"F7FF",x"FAFF",x"FCFF",x"FEFF",x"FBFF",x"FCFF",x"FCFF",x"FCFF",x"0100",x"0000",x"FFFF",x"0000",x"FEFF",x"FCFF",x"FEFF",x"FFFF",x"FEFF",x"FFFF",x"FEFF",x"0100",x"0500",x"0700",x"0A00",x"0800",x"0700",x"0400",x"0100",x"0000",x"FEFF",x"FEFF",x"F9FF",x"FBFF",x"FEFF",x"FFFF",x"FEFF",x"0200",x"0400",x"0500",x"0300",x"0200",x"0200",x"0500",x"0600",x"0600",x"0900",x"0800",x"0700",x"0700",x"0700",x"0800",x"0400",x"0400",x"0600",x"0400",x"0300",x"0100",x"0300",x"0200",x"FDFF",x"FCFF",x"FEFF",x"FEFF",x"FEFF",x"FFFF",x"FBFF",x"F9FF",x"F9FF",x"F9FF",x"FCFF",x"FAFF",x"F9FF",x"F9FF",x"FAFF",x"FDFF",x"FBFF",x"FBFF",x"FAFF",x"F8FF",x"FEFF",x"FEFF",x"FDFF",x"0400",x"0400",x"0100",x"0000",x"0100",x"0000",x"0100",x"FDFF",x"FCFF",x"FAFF",x"F9FF",x"F8FF",x"FAFF",x"FBFF",x"F9FF",x"FDFF",x"0100",x"0000",x"FCFF",x"FBFF",x"FEFF",x"FFFF",x"FEFF",x"0100",x"0400",x"0500",x"0300",x"0300",x"0200",x"0200",x"0200",x"0300",x"0600",x"0800",x"0800",x"0800",x"0600",x"0100",x"0100",x"0400",x"0500",x"0500",x"0800",x"0900",x"0900",x"0700",x"0400",x"0100",x"0100",x"0100",x"0200",x"0400",x"0300",x"0400",x"0600",x"0400",x"0100",x"0300",x"0300",x"0400",x"0300",x"0200",x"0100",x"FBFF",x"F9FF",x"FBFF",x"FDFF",x"FDFF",x"FFFF",x"FFFF",x"FEFF",x"FBFF",x"FBFF",x"FBFF",x"FFFF",x"FFFF",x"FFFF",x"0100",x"FFFF",x"FCFF",x"FBFF",x"FAFF",x"F7FF",x"FAFF",x"FEFF",x"FCFF",x"FBFF",x"FAFF",x"F8FF",x"FAFF",x"FDFF",x"0100",x"0400",x"0400",x"0100",x"0200",x"0500",x"0500",x"0600",x"0600",x"0500",x"0100",x"FFFF",x"FEFF",x"FBFF",x"FBFF",x"F9FF",x"FBFF",x"FAFF",x"F7FF",x"F6FF",x"FBFF",x"FDFF",x"FDFF",x"FBFF",x"FCFF",x"0000",x"0000",x"0100",x"0300",x"0400",x"0600",x"0700",x"0600",x"0700",x"0900",x"0900",x"0800",x"0800",x"0700",x"0300",x"0200",x"0100",x"0000",x"0100",x"0000",x"0300",x"FFFF",x"FDFF",x"0000",x"FFFF",x"FEFF",x"FDFF",x"FFFF",x"0000",x"0100",x"0500",x"0500",x"0300",x"0500",x"0100",x"0000",x"0200");	 							   
				--
				signal Zero_voice: Zero:=(x"494E", x"464F", x"4953", x"4654", x"0E00", x"0000", x"4C61", x"7666", x"3538", x"2E37", x"362E", x"3130", x"3000", x"6461", x"7461", x"BC25", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0100", x"FFFF", x"FFFF", x"0100", x"0000", x"FFFF", x"0000", x"0100", x"FFFF", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"FEFF", x"FFFF", x"FEFF", x"FEFF", x"0400", x"0600", x"0400", x"0500", x"0800", x"0400", x"0300", x"0200", x"0100", x"0100", x"FFFF", x"0200", x"0300", x"0300", x"0000", x"0000", x"0400", x"0500", x"FDFF", x"FFFF", x"FEFF", x"FDFF", x"0000", x"FEFF", x"0200", x"0300", x"0300", x"0500", x"0000", x"FEFF", x"FEFF", x"FFFF", x"0000", x"FDFF", x"FCFF", x"FAFF", x"FBFF", x"FDFF", x"FDFF", x"FBFF", x"F9FF", x"FBFF", x"FCFF", x"FBFF", x"FEFF", x"FFFF", x"FDFF", x"FFFF", x"0200", x"0000", x"0000", x"0200", x"0100", x"FEFF", x"FDFF", x"FCFF", x"FFFF", x"FFFF", x"0100", x"0900", x"0A00", x"0700", x"0400", x"0000", x"0300", x"0200", x"0000", x"0000", x"0000", x"0300", x"0000", x"FFFF", x"0400", x"0400", x"0000", x"0300", x"0600", x"0400", x"0400", x"0500", x"0100", x"0000", x"FFFF", x"0100", x"0100", x"0000", x"FFFF", x"FEFF", x"FCFF", x"FDFF", x"FDFF", x"FFFF", x"0200", x"0400", x"0300", x"0000", x"FEFF", x"FDFF", x"FBFF", x"FDFF", x"0100", x"0200", x"FFFF", x"0200", x"0000", x"FDFF", x"FDFF", x"FBFF", x"FFFF", x"0000", x"0100", x"FFFF", x"FEFF", x"FFFF", x"0100", x"0400", x"0600", x"0300", x"0000", x"FFFF", x"FFFF", x"FCFF", x"FCFF", x"FAFF", x"F8FF", x"FAFF", x"FDFF", x"FCFF", x"FEFF", x"FDFF", x"FDFF", x"0200", x"FDFF", x"FFFF", x"0000", x"FCFF", x"FBFF", x"FAFF", x"FBFF", x"FEFF", x"FDFF", x"FCFF", x"0000", x"0200", x"0100", x"0000", x"0100", x"0400", x"0800", x"0700", x"0900", x"0700", x"0200", x"0500", x"0400", x"0500", x"0700", x"0700", x"0300", x"0200", x"0600", x"0700", x"0400", x"0100", x"0300", x"0300", x"FFFF", x"FEFF", x"FFFF", x"FFFF", x"FEFF", x"FBFF", x"FDFF", x"FCFF", x"FDFF", x"FCFF", x"FEFF", x"0100", x"0300", x"0500", x"0400", x"0000", x"FFFF", x"FFFF", x"FFFF", x"0000", x"FEFF", x"F6FF", x"F4FF", x"F8FF", x"FDFF", x"FFFF", x"0000", x"0200", x"FFFF", x"0100", x"0100", x"FFFF", x"0000", x"0000", x"FEFF", x"FCFF", x"FBFF", x"FFFF", x"FEFF", x"FDFF", x"0100", x"0200", x"0200", x"0500", x"0500", x"0000", x"0200", x"0300", x"0200", x"0700", x"0300", x"0500", x"0400", x"FFFF", x"0300", x"0200", x"0000", x"FFFF", x"FFFF", x"0100", x"0200", x"0000", x"FFFF", x"FFFF", x"0200", x"0000", x"0000", x"0300", x"FEFF", x"FDFF", x"0200", x"0200", x"0100", x"0400", x"0300", x"0100", x"0100", x"0000", x"0100", x"FEFF", x"FAFF", x"FAFF", x"FDFF", x"0000", x"FEFF", x"FCFF", x"FBFF", x"FDFF", x"FEFF", x"FAFF", x"FDFF", x"FFFF", x"FAFF", x"FDFF", x"FEFF", x"FDFF", x"FDFF", x"FDFF", x"FDFF", x"FEFF", x"FFFF", x"0000", x"FFFF", x"FDFF", x"FDFF", x"FCFF", x"0200", x"0200", x"FEFF", x"0100", x"0100", x"0200", x"0600", x"0600", x"0600", x"0500", x"0500", x"0300", x"0800", x"0800", x"0500", x"0600", x"0500", x"0500", x"0600", x"0400", x"FFFF", x"0000", x"FFFF", x"FCFF", x"FCFF", x"FFFF", x"FEFF", x"FDFF", x"FBFF", x"FAFF", x"FAFF", x"FBFF", x"FBFF", x"FBFF", x"FDFF", x"FCFF", x"FBFF", x"F9FF", x"F9FF", x"FCFF", x"FFFF", x"0000", x"0600", x"0600", x"0500", x"0900", x"0800", x"0A00", x"0600", x"0200", x"0500", x"0500", x"0700", x"0600", x"0700", x"0B00", x"0B00", x"0800", x"0700", x"0600", x"0600", x"0500", x"0300", x"0200", x"0100", x"0100", x"0100", x"FDFF", x"FCFF", x"FFFF", x"F8FF", x"F8FF", x"FBFF", x"FAFF", x"F8FF", x"F5FF", x"F4FF", x"F2FF", x"F1FF", x"F3FF", x"F7FF", x"FAFF", x"0000", x"FFFF", x"FFFF", x"FBFF", x"F8FF", x"F9FF", x"FBFF", x"FBFF", x"FDFF", x"0200", x"FFFF", x"FFFF", x"FEFF", x"FDFF", x"FFFF", x"0200", x"0500", x"0400", x"0600", x"0400", x"0500", x"0A00", x"0400", x"0100", x"0100", x"0300", x"0100", x"0100", x"0000", x"0000", x"0400", x"0300", x"FEFF", x"FFFF", x"FFFF", x"0100", x"0500", x"0400", x"0300", x"0000", x"FEFF", x"FFFF", x"0000", x"0300", x"0200", x"0000", x"0200", x"0500", x"0200", x"0300", x"0700", x"0400", x"0400", x"0000", x"0200", x"0100", x"0100", x"0300", x"0200", x"0500", x"0300", x"0300", x"0200", x"FEFF", x"0100", x"FFFF", x"0100", x"0100", x"FDFF", x"0100", x"0200", x"0100", x"0000", x"FDFF", x"FFFF", x"0200", x"FEFF", x"0000", x"FEFF", x"FBFF", x"FDFF", x"FCFF", x"FDFF", x"FEFF", x"FDFF", x"FCFF", x"FBFF", x"FBFF", x"FDFF", x"FFFF", x"FEFF", x"FCFF", x"FBFF", x"0000", x"FDFF", x"FEFF", x"FCFF", x"FEFF", x"0000", x"FEFF", x"FFFF", x"0100", x"FEFF", x"FCFF", x"FCFF", x"FCFF", x"FFFF", x"FFFF", x"0200", x"0500", x"0100", x"FFFF", x"FCFF", x"FFFF", x"FFFF", x"FEFF", x"FDFF", x"0000", x"0100", x"0200", x"0200", x"0100", x"0000", x"0300", x"0500", x"0700", x"0700", x"0500", x"0200", x"0000", x"FDFF", x"FAFF", x"FAFF", x"FEFF", x"0100", x"0400", x"0400", x"0400", x"0200", x"0200", x"0800", x"0600", x"0800", x"0700", x"0600", x"0900", x"0600", x"0100", x"0000", x"0400", x"0300", x"0400", x"0200", x"0200", x"FFFF", x"FFFF", x"0100", x"0000", x"0300", x"FFFF", x"0100", x"FDFF", x"FEFF", x"FEFF", x"FCFF", x"FEFF", x"FFFF", x"FFFF", x"FEFF", x"FEFF", x"FBFF", x"F7FF", x"F8FF", x"F7FF", x"FAFF", x"FEFF", x"FCFF", x"FBFF", x"F9FF", x"FEFF", x"FBFF", x"FEFF", x"FDFF", x"FCFF", x"FEFF", x"FDFF", x"FAFF", x"FBFF", x"FCFF", x"FDFF", x"FDFF", x"0500", x"0700", x"0600", x"0100", x"0000", x"0300", x"0100", x"0100", x"FFFF", x"FFFF", x"FEFF", x"0000", x"0000", x"FFFF", x"0400", x"0300", x"0400", x"0400", x"0500", x"0600", x"0200", x"0300", x"FFFF", x"FCFF", x"FBFF", x"FBFF", x"FAFF", x"FCFF", x"0000", x"0000", x"0400", x"0200", x"0500", x"0500", x"FFFF", x"0100", x"0000", x"0300", x"0000", x"0500", x"0600", x"0400", x"0500", x"0700", x"0700", x"0300", x"0900", x"0700", x"0800", x"0300", x"0200", x"0300", x"FEFF", x"0200", x"0100", x"0200", x"0400", x"0600", x"0600", x"0100", x"FEFF", x"FBFF", x"FFFF", x"FBFF", x"FBFF", x"FEFF", x"FAFF", x"FAFF", x"F9FF", x"FCFF", x"FBFF", x"FAFF", x"FBFF", x"FBFF", x"FEFF", x"FBFF", x"FDFF", x"F9FF", x"F8FF", x"FCFF", x"FAFF", x"FAFF", x"FCFF", x"0000", x"FCFF", x"FFFF", x"0100", x"0200", x"FFFF", x"FFFF", x"0200", x"FCFF", x"0200", x"0200", x"0200", x"0200", x"0300", x"0400", x"0200", x"0000", x"0200", x"0100", x"FBFF", x"FCFF", x"F7FF", x"F5FF", x"F7FF", x"F7FF", x"FBFF", x"FBFF", x"FAFF", x"FCFF", x"FDFF", x"0100", x"0400", x"0800", x"0A00", x"0400", x"0500", x"0300", x"0400", x"0400", x"0400", x"0700", x"0900", x"0C00", x"0900", x"0A00", x"0A00", x"0400", x"0100", x"0000", x"0200", x"0200", x"FFFF", x"0000", x"0200", x"FDFF", x"FBFF", x"FEFF", x"FFFF", x"0100", x"0100", x"FFFF", x"FEFF", x"0000", x"0000", x"FFFF", x"0100", x"FDFF", x"FEFF", x"FBFF", x"FAFF", x"FCFF", x"FFFF", x"FCFF", x"FCFF", x"FCFF", x"FFFF", x"0100", x"0200", x"0100", x"0000", x"FEFF", x"FCFF", x"FCFF", x"FEFF", x"0100", x"0400", x"0100", x"0300", x"0200", x"0300", x"0000", x"0100", x"0300", x"0100", x"0500", x"0400", x"0500", x"0300", x"FDFF", x"0100", x"FDFF", x"0000", x"0000", x"FEFF", x"0000", x"FFFF", x"0200", x"0300", x"0000", x"0100", x"0200", x"0100", x"FFFF", x"FFFF", x"0300", x"0200", x"0200", x"FFFF", x"FFFF", x"FEFF", x"FFFF", x"FFFF", x"0000", x"0100", x"0200", x"0200", x"FFFF", x"0300", x"0400", x"0400", x"0500", x"FFFF", x"FCFF", x"FAFF", x"F7FF", x"F9FF", x"F7FF", x"F5FF", x"F8FF", x"FBFF", x"F9FF", x"FAFF", x"FDFF", x"FFFF", x"0100", x"FBFF", x"F7FF", x"F8FF", x"FDFF", x"FEFF", x"FFFF", x"0500", x"0600", x"0600", x"0900", x"0900", x"0600", x"0500", x"0400", x"0100", x"FFFF", x"FEFF", x"FBFF", x"FEFF", x"FFFF", x"0100", x"0600", x"0900", x"0A00", x"0E00", x"0A00", x"0C00", x"0E00", x"0900", x"0400", x"FEFF", x"0100", x"FEFF", x"FEFF", x"FEFF", x"0300", x"0400", x"0700", x"0400", x"0400", x"0300", x"FFFF", x"FFFF", x"F7FF", x"F9FF", x"F5FF", x"F4FF", x"F6FF", x"F7FF", x"FDFF", x"FDFF", x"FCFF", x"FEFF", x"0200", x"FFFF", x"FDFF", x"FAFF", x"F9FF", x"FBFF", x"F8FF", x"F8FF", x"F8FF", x"FBFF", x"FCFF", x"0200", x"FDFF", x"FAFF", x"F7FF", x"FDFF", x"0100", x"FDFF", x"0000", x"FEFF", x"FDFF", x"FFFF", x"0100", x"0400", x"0300", x"0200", x"0200", x"0200", x"0200", x"FDFF", x"F9FF", x"FBFF", x"FDFF", x"FEFF", x"FEFF", x"0200", x"0500", x"0600", x"0A00", x"0A00", x"0500", x"0600", x"0700", x"0500", x"0500", x"0400", x"0800", x"0900", x"0900", x"0B00", x"0B00", x"0B00", x"0800", x"0800", x"0700", x"0100", x"FFFF", x"FCFF", x"0400", x"0400", x"FFFF", x"0500", x"0700", x"0A00", x"0600", x"0200", x"0100", x"FFFF", x"FEFF", x"FDFF", x"0100", x"0100", x"FEFF", x"FFFF", x"0000", x"FDFF", x"FDFF", x"FFFF", x"0100", x"0300", x"FEFF", x"F6FF", x"F5FF", x"F3FF", x"F4FF", x"F5FF", x"F6FF", x"FAFF", x"F8FF", x"F5FF", x"F3FF", x"F2FF", x"F3FF", x"FDFF", x"FBFF", x"FFFF", x"FEFF", x"FDFF", x"FFFF", x"FDFF", x"FEFF", x"F8FF", x"FCFF", x"FAFF", x"F8FF", x"FEFF", x"0400", x"0500", x"0800", x"0900", x"0600", x"0900", x"0900", x"0900", x"0600", x"0600", x"0300", x"0500", x"0400", x"FEFF", x"0300", x"0400", x"0400", x"0200", x"0000", x"FDFF", x"FBFF", x"FEFF", x"FFFF", x"FFFF", x"FDFF", x"0000", x"0100", x"0400", x"0300", x"0500", x"0200", x"0200", x"0600", x"0700", x"0A00", x"0400", x"0300", x"0100", x"0300", x"0500", x"0400", x"0300", x"0000", x"FFFF", x"FDFF", x"0200", x"0200", x"0700", x"0000", x"FCFF", x"FBFF", x"F8FF", x"FBFF", x"F9FF", x"FEFF", x"FDFF", x"0000", x"0200", x"0300", x"0600", x"0100", x"0000", x"0000", x"0200", x"0000", x"0700", x"0800", x"0700", x"0300", x"0000", x"0100", x"FDFF", x"0000", x"FFFF", x"0300", x"FFFF", x"FDFF", x"FBFF", x"FAFF", x"FDFF", x"FFFF", x"FDFF", x"FFFF", x"FFFF", x"0000", x"FEFF", x"FBFF", x"FCFF", x"FAFF", x"FAFF", x"FBFF", x"FBFF", x"F9FF", x"F9FF", x"FEFF", x"0200", x"0200", x"FAFF", x"FAFF", x"F8FF", x"FBFF", x"0000", x"0300", x"0700", x"0A00", x"0900", x"0700", x"0500", x"0500", x"0400", x"0200", x"0200", x"0100", x"0100", x"0100", x"FEFF", x"0200", x"0200", x"0500", x"0100", x"FFFF", x"FCFF", x"F8FF", x"FAFF", x"FAFF", x"FFFF", x"FDFF", x"0000", x"0500", x"0600", x"0700", x"0600", x"0500", x"0200", x"FEFF", x"FDFF", x"0300", x"FEFF", x"FCFF", x"F7FF", x"F7FF", x"F8FF", x"F6FF", x"F6FF", x"F8FF", x"FAFF", x"FFFF", x"FFFF", x"0000", x"0000", x"0500", x"0A00", x"0900", x"0600", x"0500", x"0300", x"FFFF", x"0200", x"0500", x"0400", x"0300", x"0200", x"0300", x"0600", x"0300", x"0700", x"0300", x"0100", x"0600", x"0200", x"FFFF", x"FEFF", x"FEFF", x"0000", x"FEFF", x"FDFF", x"FFFF", x"FFFF", x"FFFF", x"FEFF", x"FFFF", x"0000", x"0100", x"0200", x"0100", x"0100", x"0000", x"0100", x"0000", x"FEFF", x"FDFF", x"FCFF", x"FDFF", x"FEFF", x"FDFF", x"FCFF", x"F8FF", x"FDFF", x"FDFF", x"FCFF", x"0000", x"0300", x"0300", x"0300", x"0100", x"0000", x"FEFF", x"0300", x"0200", x"0100", x"FFFF", x"FEFF", x"0200", x"0100", x"0300", x"0100", x"0100", x"0200", x"FBFF", x"F8FF", x"FAFF", x"FBFF", x"FBFF", x"0200", x"0400", x"0600", x"0600", x"0500", x"0300", x"0000", x"0100", x"FEFF", x"0100", x"FFFF", x"FFFF", x"0300", x"FFFF", x"0200", x"0600", x"0200", x"0000", x"FFFF", x"0100", x"FEFF", x"F9FF", x"F7FF", x"F8FF", x"F6FF", x"F9FF", x"FEFF", x"FBFF", x"FEFF", x"0000", x"F9FF", x"F9FF", x"FAFF", x"FBFF", x"0200", x"0100", x"0300", x"0500", x"0500", x"0300", x"0600", x"0800", x"0900", x"0A00", x"0700", x"0400", x"0300", x"0000", x"FCFF", x"FBFF", x"FEFF", x"0200", x"0400", x"0700", x"0400", x"0200", x"FFFF", x"FBFF", x"FBFF", x"FFFF", x"0300", x"0300", x"0100", x"FFFF", x"FFFF", x"FDFF", x"FCFF", x"FFFF", x"FEFF", x"0300", x"FEFF", x"FCFF", x"FFFF", x"FFFF", x"0200", x"0600", x"0400", x"0400", x"0300", x"FCFF", x"0400", x"0500", x"0300", x"0200", x"FFFF", x"FFFF", x"FBFF", x"FEFF", x"FAFF", x"FDFF", x"0200", x"0100", x"FEFF", x"0300", x"0300", x"0000", x"0500", x"0400", x"0300", x"0400", x"FEFF", x"FDFF", x"FCFF", x"F9FF", x"FFFF", x"FFFF", x"FEFF", x"0100", x"0300", x"0300", x"0300", x"FEFF", x"FBFF", x"FDFF", x"FFFF", x"FFFF", x"0100", x"0000", x"FFFF", x"FBFF", x"FAFF", x"FDFF", x"FDFF", x"FBFF", x"FBFF", x"FFFF", x"0100", x"0400", x"0500", x"0600", x"0000", x"0200", x"0100", x"0300", x"0500", x"0400", x"0500", x"0600", x"0500", x"0100", x"0000", x"FFFF", x"FCFF", x"FDFF", x"0000", x"0300", x"0700", x"0300", x"0300", x"0300", x"FDFF", x"FEFF", x"FEFF", x"F9FF", x"FAFF", x"F9FF", x"FBFF", x"FFFF", x"0100", x"0100", x"0100", x"0500", x"0200", x"0400", x"0500", x"0600", x"0100", x"0000", x"0400", x"0000", x"0100", x"0300", x"0300", x"0500", x"0200", x"0400", x"FFFF", x"FCFF", x"FAFF", x"F9FF", x"F8FF", x"FCFF", x"FCFF", x"FAFF", x"F9FF", x"FFFF", x"FFFF", x"FAFF", x"FBFF", x"FBFF", x"FAFF", x"FAFF", x"FAFF", x"F6FF", x"F6FF", x"F6FF", x"FBFF", x"FAFF", x"FEFF", x"FDFF", x"FFFF", x"0200", x"0100", x"0100", x"0000", x"FFFF", x"0300", x"0300", x"0300", x"0300", x"0000", x"FDFF", x"FEFF", x"0000", x"0000", x"0100", x"0600", x"0A00", x"0A00", x"0B00", x"1000", x"0F00", x"0D00", x"0B00", x"0A00", x"0C00", x"0E00", x"0E00", x"0800", x"FFFF", x"F9FF", x"F8FF", x"F8FF", x"FBFF", x"FDFF", x"FAFF", x"FAFF", x"FBFF", x"FEFF", x"FDFF", x"FCFF", x"FEFF", x"0100", x"0400", x"0300", x"0500", x"0400", x"0000", x"0100", x"FDFF", x"FEFF", x"FFFF", x"FEFF", x"0000", x"0200", x"0100", x"FFFF", x"0000", x"0400", x"0200", x"0300", x"0100", x"FEFF", x"FDFF", x"FBFF", x"FBFF", x"FBFF", x"F6FF", x"F4FF", x"F8FF", x"FBFF", x"FAFF", x"0100", x"0400", x"0500", x"0200", x"0400", x"0100", x"FCFF", x"FBFF", x"FCFF", x"FBFF", x"FDFF", x"FCFF", x"FAFF", x"FDFF", x"FBFF", x"FEFF", x"0100", x"0200", x"0500", x"0300", x"0100", x"0000", x"0100", x"0400", x"0000", x"0100", x"0200", x"0200", x"FDFF", x"FBFF", x"FAFF", x"FEFF", x"0200", x"0300", x"FFFF", x"0100", x"0300", x"0300", x"0000", x"FCFF", x"0000", x"0000", x"FFFF", x"0200", x"0300", x"0000", x"FFFF", x"0200", x"0500", x"0B00", x"0800", x"0700", x"0700", x"0300", x"0600", x"0700", x"0300", x"0300", x"0500", x"0500", x"0500", x"0000", x"FEFF", x"FCFF", x"FBFF", x"FBFF", x"FEFF", x"0100", x"0300", x"0600", x"0100", x"0300", x"0200", x"0000", x"0100", x"FEFF", x"FFFF", x"FFFF", x"FCFF", x"FCFF", x"FDFF", x"F9FF", x"FBFF", x"F8FF", x"FAFF", x"FCFF", x"FBFF", x"FFFF", x"0100", x"0100", x"0100", x"0500", x"0300", x"0300", x"0000", x"FCFF", x"FBFF", x"FDFF", x"0100", x"0000", x"0100", x"0200", x"FFFF", x"0000", x"0000", x"FFFF", x"FEFF", x"FFFF", x"0400", x"0300", x"0400", x"0200", x"0000", x"0100", x"FEFF", x"FDFF", x"FEFF", x"FBFF", x"FBFF", x"FEFF", x"FAFF", x"FCFF", x"FEFF", x"FFFF", x"FDFF", x"FBFF", x"FEFF", x"0100", x"0200", x"FFFF", x"0300", x"0200", x"0000", x"0200", x"FCFF", x"0200", x"0300", x"0200", x"0100", x"0000", x"FEFF", x"FDFF", x"0400", x"0800", x"0900", x"0600", x"0400", x"0700", x"0400", x"0800", x"0700", x"0900", x"0900", x"0600", x"0600", x"0600", x"0600", x"0600", x"0500", x"FDFF", x"FBFF", x"F8FF", x"F7FF", x"F8FF", x"F8FF", x"FAFF", x"F9FF", x"F7FF", x"F9FF", x"FBFF", x"FFFF", x"0400", x"0200", x"FEFF", x"FDFF", x"FEFF", x"FBFF", x"F8FF", x"FCFF", x"FDFF", x"FDFF", x"0300", x"0200", x"0200", x"0300", x"0100", x"0300", x"FFFF", x"FDFF", x"0200", x"0100", x"FEFF", x"FBFF", x"F8FF", x"F9FF", x"FAFF", x"FDFF", x"FDFF", x"FDFF", x"FAFF", x"FCFF", x"FFFF", x"FCFF", x"0100", x"0300", x"0600", x"0700", x"0300", x"0400", x"0400", x"0300", x"0300", x"0300", x"0100", x"0100", x"0300", x"0500", x"0100", x"0200", x"0300", x"FBFF", x"FFFF", x"FFFF", x"FBFF", x"FBFF", x"FAFF", x"FDFF", x"0000", x"0200", x"0000", x"0400", x"0500", x"0200", x"0100", x"FDFF", x"F8FF", x"F8FF", x"FBFF", x"FEFF", x"0000", x"0300", x"0700", x"0600", x"0900", x"0A00", x"0B00", x"0800", x"0800", x"0300", x"0200", x"0400", x"FFFF", x"FBFF", x"FCFF", x"FEFF", x"FFFF", x"0100", x"0400", x"0500", x"0600", x"0500", x"0400", x"0700", x"0600", x"0300", x"0200", x"FEFF", x"FCFF", x"FAFF", x"F9FF", x"F9FF", x"F6FF", x"F7FF", x"F7FF", x"F9FF", x"F8FF", x"FBFF", x"FEFF", x"FFFF", x"0400", x"0400", x"0400", x"0400", x"0700", x"0700", x"0000", x"FEFF", x"FDFF", x"FAFF", x"0100", x"FFFF", x"FFFF", x"0500", x"0800", x"0700", x"0400", x"0200", x"FEFF", x"FEFF", x"FDFF", x"F9FF", x"FDFF", x"FDFF", x"0000", x"FFFF", x"0200", x"0100", x"FDFF", x"0300", x"FFFF", x"0800", x"0400", x"0700", x"1600", x"0E00", x"2700", x"1400", x"1800", x"FEFF", x"EEFF", x"DCFF", x"CEFF", x"D3FF", x"CBFF", x"DBFF", x"E0FF", x"ECFF", x"FDFF", x"0400", x"2100", x"1F00", x"3900", x"3C00", x"3100", x"3A00", x"1D00", x"2100", x"0300", x"EFFF", x"DAFF", x"C3FF", x"B8FF", x"ADFF", x"B1FF", x"B9FF", x"D6FF", x"DDFF", x"EAFF", x"EDFF", x"EDFF", x"EFFF", x"F5FF", x"FDFF", x"0600", x"1000", x"1900", x"1F00", x"2600", x"3800", x"3F00", x"5400", x"5900", x"6A00", x"6F00", x"6A00", x"5B00", x"4900", x"2F00", x"1500", x"F5FF", x"DFFF", x"C2FF", x"BBFF", x"A7FF", x"A0FF", x"9CFF", x"9BFF", x"A3FF", x"B1FF", x"C1FF", x"DCFF", x"F7FF", x"1000", x"3400", x"4200", x"5A00", x"6300", x"6C00", x"6F00", x"6800", x"5F00", x"5400", x"2D00", x"1900", x"EEFF", x"CAFF", x"A0FF", x"80FF", x"63FF", x"4DFF", x"47FF", x"48FF", x"53FF", x"70FF", x"86FF", x"A2FF", x"B5FF", x"C8FF", x"D6FF", x"EDFF", x"0300", x"2E00", x"5D00", x"9F00", x"E400", x"2801", x"6C01", x"9B01", x"A601", x"8B01", x"4101", x"DA00", x"4F00", x"C8FF", x"4AFF", x"E2FE", x"90FE", x"5FFE", x"45FE", x"4DFE", x"45FE", x"6DFE", x"6EFE", x"ABFE", x"C6FE", x"17FF", x"4DFF", x"B2FF", x"0600", x"7F00", x"FD00", x"BF01", x"8202", x"7003", x"2B04", x"B604", x"AE04", x"3304", x"2E03", x"DA01", x"6100", x"DAFE", x"9BFD", x"94FC", x"E2FB", x"80FB", x"56FB", x"86FB", x"FDFB", x"99FC", x"7EFD", x"72FE", x"47FF", x"ECFF", x"4700", x"5000", x"3800", x"0100", x"F4FF", x"4700", x"1601", x"3902", x"9A03", x"9604", x"5105", x"1C05", x"8104", x"3E03", x"2402", x"E000", x"1C00", x"59FF", x"FAFE", x"6EFE", x"FDFD", x"53FD", x"A6FC", x"35FC", x"F4FB", x"0DFC", x"80FC", x"EDFC", x"7CFD", x"ECFD", x"41FE", x"71FE", x"72FE", x"7DFE", x"94FE", x"EBFE", x"68FF", x"9300", x"F601", x"C303", x"7205", x"A506", x"0407", x"9206", x"6305", x"E503", x"8902", x"7401", x"C400", x"5000", x"D3FF", x"40FF", x"96FE", x"ACFD", x"E7FC", x"3DFC", x"9EFB", x"67FB", x"6FFB", x"B0FB", x"08FC", x"6FFC", x"E4FC", x"4DFD", x"ADFD", x"06FE", x"5EFE", x"B8FE", x"36FF", x"1800", x"A101", x"7403", x"DA05", x"9907", x"E108", x"D108", x"0008", x"4606", x"A204", x"0803", x"0202", x"FF00", x"4000", x"59FF", x"4FFE", x"0BFD", x"F2FB", x"F0FA", x"2AFA", x"3DFA", x"3EFA", x"8DFA", x"19FB", x"9AFB", x"25FC", x"A1FC", x"20FD", x"65FD", x"C6FD", x"FCFD", x"71FE", x"08FF", x"6400", x"2502", x"6D04", x"EC06", x"EF08", x"3A0A", x"5B0A", x"7509", x"C007", x"D705", x"EE03", x"9002", x"4201", x"5900", x"20FF", x"B0FD", x"05FC", x"8CFA", x"12F9", x"78F8", x"10F8", x"45F8", x"BEF8", x"9CF9", x"30FA", x"1EFB", x"D4FB", x"79FC", x"21FD", x"87FD", x"11FE", x"6CFE", x"27FF", x"EF00", x"0703", x"E605", x"A908", x"7D0A", x"560B", x"EB0A", x"8A09", x"0308", x"7306", x"3A05", x"F903", x"A402", x"E000", x"17FF", x"1CFD", x"69FB", x"24F9", x"19F8", x"14F7", x"51F7", x"07F8", x"4AF9", x"7CFA", x"7DFB", x"20FC", x"57FC", x"87FC", x"31FD", x"0DFD", x"F9FD", x"57FE", x"6C00", x"8802", x"EB05", x"1709", x"B80B", x"290D", x"E50C", x"6C0B", x"3809", x"2607", x"BD04", x"2D03", x"9701", x"EDFF", x"EFFD", x"4FFC", x"62FA", x"14F8", x"4EF7", x"60F6", x"29F6", x"69F7", x"2DF8", x"D8F9", x"C6FA", x"1BFC", x"2AFC", x"A7FC", x"97FC", x"84FC", x"DCFC", x"7DFD", x"2400", x"A402", x"F406", x"9F0A", x"B30D", x"330F", x"890E", x"A00C", x"9509", x"F406", x"3804", x"C002", x"2B01", x"D0FF", x"5EFE", x"88FC", x"8CFA", x"B9F8", x"68F7", x"97F6", x"E1F6", x"38F7", x"FDF7", x"73F8", x"A3F8", x"62F9", x"2AFA", x"70FA", x"0AFB", x"6BFB", x"64FB", x"D6FC", x"69FF", x"B702", x"9008", x"AD0C", x"0911", x"5112", x"7911", x"A90E", x"B90A", x"3D07", x"5104", x"9002", x"2001", x"3100", x"DDFE", x"27FD", x"14FB", x"E2F8", x"0EF7", x"A6F5", x"33F5", x"6BF5", x"B2F5", x"0DF7", x"7FF7", x"17F9", x"FFF8", x"5CF9", x"13F8", x"79F9", x"D5F8", x"AAFC", x"3100", x"A306", x"640D", x"B112", x"5616", x"BF15", x"6713", x"A10E", x"A409", x"F005", x"6403", x"6B01", x"EE00", x"CCFE", x"DAFC", x"B9F9", x"D3F7", x"50F5", x"D8F4", x"0EF5", x"34F5", x"26F6", x"8CF6", x"D6F6", x"1DF8", x"FDF7", x"EEF8", x"36F8", x"FFF8", x"A3F7", x"97FB", x"23FF", x"D406", x"D40E", x"3015", x"C219", x"0619", x"E215", x"620F", x"6A0A", x"8F04", x"AE02", x"0B01", x"DCFF", x"F0FE", x"02FC", x"4FF9", x"70F7", x"CFF4", x"62F3", x"D5F2", x"10F3", x"3DF4", x"25F6", x"3DF7", x"38F8", x"13F8", x"6DF8", x"6EF6", x"CFF6", x"EBF4", x"B7FB", x"28FF", x"470A", x"E911", x"791A", x"941D", x"2D1C", x"2C16", x"C20D", x"8606", x"BB00", x"C9FE", x"07FE", x"3DFF", x"35FE", x"6EFD", x"75F9", x"D0F6", x"F3F3", x"3FF2", x"A4F3", x"48F5", x"F9F6", x"00F8", x"87F8", x"52F7", x"7FF6", x"48F4", x"39F4", x"B4F1", x"89F7", x"59FD", x"4808", x"2B13", x"761B", x"4020", x"4A1E", x"FF18", x"770E", x"6A07", x"AEFF", x"24FE", x"5EFC", x"33FF", x"F7FE", x"A5FD", x"5FFA", x"14F8", x"5EF4", x"0EF3", x"52F4", x"C9F6", x"02F7", x"F0F9", x"FAF8", x"9FF6", x"75F5", x"8BF0", x"3DF0", x"49ED", x"97F8", x"A4FC", x"460F", x"8018", x"3D24", x"B524", x"9721", x"3F17", x"D00B", x"A501", x"EDFA", x"18FA", x"82FA", x"E0FD", x"0BFD", x"B3FB", x"E0F8", x"45F5", x"DEF1", x"8FF2", x"A2F4", x"A9F8", x"B0F9", x"61FC", x"B0FA", x"25F8", x"72F5", x"ECEF", x"9CE7", x"A1F3", x"08F7", x"280E", x"4319", x"562A", x"0B2C", x"5529", x"701B", x"8A0B", x"6AFD", x"F4F3", x"78F0", x"BCF1", x"8AF6", x"ADFA", x"0AFC", x"F3F8", x"94F5", x"FFF2", x"9BF0", x"A4F2", x"13F5", x"6DF8", x"7BFA", x"9EF9", x"ADF5", x"54F4", x"DCEA", x"F9F3", x"D3FB", x"890E", x"3023", x"022E", x"4837", x"232C", x"1A1E", x"0305", x"9EF6", x"C1E8", x"68EB", x"DAEC", x"D2F7", x"87FB", x"60FF", x"04FC", x"1AF7", x"EAEE", x"F9ED", x"09F0", x"BDF4", x"D5FA", x"C6FC", x"96FB", x"A1F7", x"F7F0", x"16EA", x"BDFC", x"0A01", x"D222", x"792B", x"9D3E", x"1F35", x"332A", x"510B", x"18F5", x"69E3", x"A8E0", x"DCE6", x"B8F2", x"D1FB", x"A700", x"66FC", x"A9F4", x"7EEC", x"3AE9", x"8EEA", x"D6F0", x"78F8", x"B8FD", x"37FE", x"D5F7", x"82F3", x"24E8", x"FBFF", x"E904", x"2B2F", x"0E38", x"104E", x"D33E", x"AB2C", x"7107", x"67EB", x"40D8", x"E5D5", x"C6E0", x"51F0", x"EEFE", x"CE03", x"A9FD", x"04F3", x"C1E6", x"80E2", x"5FE3", x"27EC", x"E4F3", x"5EFE", x"CCF9", x"20FC", x"92E9", x"49F2", x"7F00", x"2812", x"6C3B", x"3F42", x"9058", x"983B", x"352B", x"4DF8", x"31E5", x"4FCE", x"04DA", x"30E4", x"4AFC", x"F905", x"3B09", x"C4FC", x"43EC", x"F7DF", x"ADDA", x"87E0", x"30EA", x"1EF6", x"EDF7", x"14FC", x"95ED", x"D3E9", x"7300", x"8F04", x"F935", x"323B", x"5758", x"2E45", x"6334", x"1F0B", x"C3EB", x"1DD7", x"5BD5", x"27E3", x"D9F5", x"D407", x"4809", x"3503", x"77EE", x"99E2", x"DAD9", x"93DF", x"14E4", x"36F5", x"02F6", x"52FD", x"C1EF", x"7EE6", x"29FF", x"C5FF", x"8D30", x"CB37", x"E551", x"9F45", x"5B30", x"DE0D", x"56E8", x"C6D9", x"73D8", x"42EC", x"9EFF", x"6D11", x"AB0F", x"A904", x"E2EB", x"5DDC", x"DAD2", x"0BD9", x"65E2", x"ADF5", x"03F9", x"97FD", x"8FF2", x"AEE3", x"E202", x"5AFD", x"7D34", x"0337", x"1352", x"4C41", x"F729", x"EA08", x"34E3", x"88D5", x"76D5", x"73EE", x"7B01", x"BC1A", x"B713", x"6A0D", x"38EF", x"D6DF", x"17CF", x"CAD7", x"08E2", x"57F4", x"59FE", x"AAFC", x"3DFB", x"3EE2", x"A003", x"3BF9", x"A127", x"2334", x"5F43", x"0945", x"F525", x"8E13", x"26E5", x"B5DD", x"D6CD", x"3DEA", x"8BF7", x"AF16", x"1418", x"4212", x"4800", x"26E8", x"09E1", x"ABD5", x"94E7", x"84EA", x"E2FF", x"6AF8", x"22FF", x"A1E8", x"23EA", x"57FB", x"9BFA", x"542D", x"322A", x"B549", x"9737", x"6727", x"460A", x"7DE6", x"9BE1", x"4CD3", x"2AF0", x"B9F9", x"AE11", x"910F", x"DE07", x"7BFA", x"7DE9", x"7FEB", x"AAE4", x"48F7", x"BDF6", x"EB03", x"0BFB", x"69FA", x"B0E9", x"F6E1", x"09F5", x"A5F0", x"BD1D", x"0622", x"053C", x"1A39", x"3F26", x"A016", x"BBF1", x"F4ED", x"32DF", x"71EB", x"BDF7", x"6D00", x"F10B", x"F2FF", x"9400", x"E6F1", x"FEF4", x"9DF0", x"88F8", x"6AFE", x"08FD", x"E400", x"18F2", x"66F4", x"DADD", x"3DE9", x"5AF2", x"D9FB", x"4721", x"B423", x"083B", x"762C", x"A31F", x"760B", x"00F4", x"BFF0", x"E4E6", x"2DF0", x"9BF9", x"8F00", x"3105", x"D6FF", x"C2FD", x"32F8", x"C0F9", x"B5F8", x"72FA", x"B1FB", x"3BFA", x"DBF8", x"7EEE", x"9DEE", x"46DE", x"65E9", x"95F8", x"3302", x"C226", x"D726", x"8239", x"B629", x"A519", x"1607", x"EFEE", x"2AEB", x"5AE5", x"84ED", x"7AF9", x"AD06", x"2B0B", x"130A", x"FF04", x"D2FC", x"22FB", x"54F5", x"F8F4", x"6BF5", x"9DF3", x"81F5", x"A9EB", x"F1ED", x"E5DE", x"16E8", x"C801", x"6E05", x"0231", x"142F", x"E03B", x"FA2B", x"780F", x"57FE", x"D1E0", x"4FE1", x"DFE0", x"F9EB", x"5202", x"F512", x"BB18", x"A913", x"3206", x"6BF6", x"C0F1", x"74EC", x"6DEF", x"84F4", x"DCF5", x"58F6", x"25E9", x"02E8", x"BFD0", x"A7F1", x"3C05", x"961C", x"404A", x"9F3A", x"FC43", x"591A", x"3FF9", x"ABE2", x"4FCE", x"CFD9", x"D6EC", x"00FD", x"EE1E", x"E921", x"AE19", x"DB0B", x"8AEE", x"90EB", x"2FE5", x"1CEC", x"04F7", x"A6F8", x"89FA", x"03E9", x"C1E0", x"75CE", x"8FDB", x"E114", x"9E18", x"255E", x"494E", x"AB3D", x"8326", x"B0E2", x"BBD5", x"FFCA", x"73CE", x"3C01", x"F608", x"F32E", x"AA2A", x"8D0A", x"F4FF", x"7ED9", x"6DE1", x"7BE6", x"24EF", x"E204", x"4CFD", x"7DFA", x"A2E1", x"A0D7", x"31BF", x"70FB", x"501A", x"933A", x"8A6D", x"2C40", x"A431", x"E501", x"8FC7", x"15D0", x"EBCE", x"C1EA", x"9C1C", x"6220", x"4034", x"5E14", x"4BF2", x"E0E1", x"B0D0", x"1DE6", x"70F4", x"2C04", x"B90B", x"F4FB", x"0BE4", x"C1D4", x"E9BC", x"EEDD", x"422A", x"6B31", x"9C6D", x"CD53", x"951D", x"E804", x"0ACC", x"F1BE", x"B2E7", x"97F5", x"C51F", x"D433", x"9820", x"D30A", x"C2EA", x"BED2", x"19DC", x"7BEB", x"44FD", x"CE0A", x"6B04", x"47F7", x"4CDB", x"E0CC", x"53C2", x"05DA", x"D638", x"A63F", x"6F60", x"A156", x"900B", x"ACED", x"17D3", x"40C1", x"E6F6", x"A519", x"5924", x"1A30", x"F015", x"97EA", x"ECE1", x"5DD5", x"EFE0", x"3801", x"380A", x"100B", x"7205", x"85EC", x"78D6", x"1CCB", x"D0CF", x"73D3", x"3B32", x"5751", x"FE46", x"BB4E", x"4410", x"80D9", x"C3DA", x"ABD5", x"F1F1", x"A025", x"A52D", x"291B", x"FB0E", x"89EE", x"05D7", x"7FE3", x"CDED", x"EAFA", x"8F12", x"880B", x"E3FB", x"8CF2", x"11E1", x"25CC", x"30D8", x"B4D6", x"9803", x"9853", x"614A", x"953D", x"B129", x"09EE", x"33CE", x"76DD", x"D0F0", x"910E", x"792B", x"AA24", x"E204", x"BCF6", x"62E7", x"C9DB", x"80ED", x"9FFD", x"0305", x"AF0C", x"3A07", x"EDF4", x"98EB", x"6AE2", x"B2D2", x"39D9", x"67DF", x"671C", x"7E50", x"B345", x"EF33", x"2B15", x"69E4", x"D9CF", x"FBE0", x"3602", x"BC19", x"2329", x"AF1D", x"7EF9", x"76EB", x"20E6", x"46E3", x"03F5", x"C207", x"970C", x"6F0B", x"9904", x"0DF8", x"A9E8", x"91E2", x"6FD9", x"6CDA", x"A9DF", x"D703", x"EF42", x"DC48", x"4B31", x"F61B", x"BFF9", x"CFD3", x"2FD6", x"3FFA", x"AB16", x"0B21", x"061F", x"3404", x"02EA", x"0AE6", x"F6E7", x"BFF2", x"8E05", x"8D13", x"1113", x"DB09", x"B1FE", x"78EE", x"52E0", x"8CDC", x"49DA", x"65DF", x"5BE2", x"1117", x"5C4B", x"4E43", x"882A", x"2410", x"1DEE", x"2ED3", x"4CDC", x"9604", x"8A20", x"921C", x"9E10", x"03FE", x"95DF", x"76DD", x"7EF4", x"8903", x"F00F", x"011B", x"D113", x"0502", x"E6F2", x"D3E9", x"9DDF", x"9FE2", x"7DE9", x"A5E9", x"EAE7", x"F7F5", x"632D", x"E549", x"2133", x"5C18", x"0007", x"DCE7", x"89D1", x"A6E4", x"FA0C", x"421D", x"0717", x"7E0B", x"4BF5", x"C1E2", x"5AE8", x"2000", x"D20E", x"D010", x"4210", x"9B07", x"13F8", x"44EE", x"46ED", x"38EA", x"4EE8", x"BAEC", x"8BEB", x"08E8", x"C5EF", x"E71D", x"3246", x"0F3D", x"E61B", x"7502", x"5AE9", x"85D5", x"78DC", x"7203", x"3F25", x"B623", x"D60C", x"4FF9", x"9FE7", x"39E0", x"4BF2", x"EF0B", x"9E16", x"BC12", x"6D0C", x"4B02", x"F8F4", x"4FED", x"59E8", x"DAE8", x"DBEF", x"CBF7", x"0EF8", x"7EF4", x"EFEE", x"050A", x"202B", x"772B", x"A418", x"FD07", x"7CFB", x"2CEE", x"50E9", x"CAFA", x"D414", x"C819", x"2006", x"BFF3", x"B7ED", x"E2EC", x"88F8", x"2A0C", x"9F16", x"5511", x"8404", x"18F9", x"33F3", x"1CF4", x"CCF9", x"BAFD", x"CDFC", x"79F9", x"38EF", x"81E1", x"E2DA", x"23E6", x"7713", x"363C", x"4F3D", x"1B22", x"CE02", x"C2EA", x"83DD", x"0AE0", x"D7FA", x"661A", x"651F", x"550E", x"D8FB", x"ABF0", x"C2EC", x"30F4", x"DE01", x"360D", x"2010", x"120B", x"4B08", x"E605", x"FAFC", x"40F3", x"36ED", x"71EC", x"DBED", x"52EF", x"91EF", x"5FF1", x"AFF2", x"0805", x"AC24", x"0731", x"4E1E", x"6205", x"63FA", x"56F2", x"9EEB", x"36F4", x"9109", x"5614", x"FE0B", x"1DFC", x"DDF3", x"66F3", x"85F6", x"C300", x"2B0F", x"CE14", x"940F", x"E708", x"9700", x"42F6", x"79F0", x"73EF", x"BAEF", x"A1F3", x"52F5", x"81F2", x"54EF", x"1DEF", x"F8F0", x"BD03", x"EF23", x"B731", x"C523", x"8C09", x"02F8", x"54F0", x"ECEC", x"9EF1", x"9B01", x"590F", x"4C0D", x"9C01", x"A6F8", x"8CF6", x"FAFA", x"2B05", x"5010", x"8614", x"E10C", x"96FF", x"D2F8", x"94F4", x"D9EE", x"EEEE", x"67F4", x"C1F9", x"DDFB", x"7CF7", x"C4F3", x"1EF5", x"D8F9", x"0BFA", x"BAFF", x"E213", x"B321", x"951B", x"CE08", x"ABFB", x"2FF8", x"1FF7", x"7AF7", x"10FF", x"3E0A", x"6E0D", x"5908", x"1002", x"6700", x"0203", x"7704", x"7103", x"2D01", x"B7FC", x"C2FA", x"E5FA", x"66F9", x"99F7", x"E1F7", x"40F8", x"9CF8", x"B6F8", x"86F7", x"39F7", x"06F9", x"4BFA", x"ABFB", x"3FFC", x"ECFD", x"0809", x"1615", x"0C15", x"1B0C", x"6E07", x"1B07", x"AF04", x"5C00", x"65FF", x"B802", x"1605", x"2B03", x"4001", x"5600", x"4BFF", x"A4FE", x"79FE", x"5BFE", x"60FD", x"84FC", x"1BFD", x"97FD", x"40FB", x"F4F7", x"00F6", x"BDF5", x"8CF6", x"9CF6", x"A3F7", x"EBFA", x"1FFE", x"19FE", x"9FFB", x"C4FB", x"DCFE", x"B106", x"B612", x"2F19", x"7815", x"750D", x"2806", x"E700", x"44FE", x"09FF", x"3702", x"B503", x"5E02", x"9100", x"2EFF", x"82FB", x"6CF8", x"BEF9", x"7FFD", x"7CFF", x"54FE", x"61FC", x"61FA", x"19F8", x"CBF6", x"AAF8", x"06FB", x"48FB", x"FEFA", x"83FA", x"5FFA", x"C8FC", x"6F01", x"6005", x"7A06", x"D605", x"8905", x"DB06", x"CE08", x"390B", x"4A0C", x"D109", x"BF05", x"B403", x"E402", x"2A01", x"43FF", x"FCFE", x"2AFE", x"39FC", x"DFFA", x"E3FA", x"E6FA", x"92F9", x"D0F8", x"11FA", x"80FB", x"ECFB", x"20FD", x"8AFE", x"FEFD", x"A4FC", x"3CFD", x"9FFE", x"F9FE", x"ADFF", x"1702", x"3204", x"4903", x"4301", x"4401", x"8601", x"FF00", x"CC02", x"6607", x"BA0A", x"8F09", x"6805", x"FB01", x"2D00", x"39FF", x"25FF", x"26FF", x"12FF", x"47FE", x"55FC", x"78FA", x"D8F9", x"EBFA", x"59FC", x"AFFD", x"35FF", x"96FF", x"F9FE", x"B8FE", x"37FF", x"4BFF", x"13FF", x"A0FF", x"D6FF", x"5BFF", x"0EFF", x"6FFF", x"A4FF", x"3000", x"4C02", x"AB04", x"4E05", x"1704", x"5F03", x"3004", x"7903", x"4C01", x"0700", x"F1FF", x"C4FF", x"33FE", x"22FD", x"55FD", x"4DFD", x"95FD", x"16FF", x"4700", x"F7FF", x"C7FF", x"EEFF", x"76FF", x"93FE", x"6CFE", x"CCFE", x"E6FE", x"CBFE", x"72FF", x"5300", x"6600", x"2700", x"8300", x"FB00", x"FD00", x"B700", x"6A00", x"5101", x"DF02", x"5002", x"0901", x"1901", x"CC00", x"21FF", x"0BFE", x"66FE", x"98FE", x"4FFE", x"E1FE", x"8DFF", x"4F00", x"3901", x"A100", x"92FF", x"90FF", x"87FF", x"6BFF", x"F6FE", x"5CFF", x"6300", x"D900", x"EE00", x"8800", x"3300", x"ED00", x"0E02", x"6802", x"B701", x"9E00", x"75FF", x"16FE", x"74FD", x"FCFD", x"A9FF", x"4301", x"A901", x"2001", x"0600", x"A9FE", x"D8FD", x"2DFE", x"2DFF", x"A2FF", x"B6FF", x"92FF", x"86FF", x"C3FE", x"FAFE", x"5A00", x"EC00", x"1701", x"2402", x"E402", x"6001", x"BCFF", x"8FFF", x"A1FF", x"79FF", x"5500", x"3F01", x"F700", x"4A00", x"F1FF", x"9FFF", x"23FF", x"96FF", x"D400", x"1A01", x"2400", x"8EFF", x"B7FF", x"DAFE", x"B6FD", x"EFFD", x"DFFE", x"32FF", x"FCFE", x"6AFF", x"C9FF", x"6BFF", x"E6FF", x"3801", x"9A01", x"C300", x"9100", x"C300", x"8700", x"AC00", x"4101", x"4701", x"9100", x"0900", x"B0FF", x"8DFF", x"A2FF", x"2600", x"7100", x"1D00", x"2F00", x"8500", x"2000", x"6CFF", x"15FF", x"7CFF", x"C0FF", x"75FF", x"64FF", x"B1FF", x"D1FF", x"ABFF", x"3BFF", x"0FFF", x"1AFF", x"D7FF", x"A100", x"3100", x"1C00", x"0101", x"7E01", x"7B01", x"6F01", x"3401", x"6B00", x"1000", x"AD00", x"D100", x"AFFF", x"C0FE", x"F1FE", x"33FF", x"21FF", x"82FF", x"2300", x"ECFF", x"BEFF", x"7EFF", x"2BFF", x"43FF", x"DBFF", x"3700", x"F1FF", x"0400", x"F6FF", x"52FF", x"2AFF", x"9FFF", x"4900", x"7000", x"B500", x"3601", x"EE00", x"7D00", x"8400", x"BD00", x"7700", x"6E00", x"E800", x"9500", x"F3FF", x"FDFF", x"1F00", x"9DFF", x"1EFF", x"61FF", x"7DFF", x"1FFF", x"69FF", x"EEFF", x"C6FF", x"3EFF", x"28FF", x"51FF", x"8DFF", x"0C00", x"2100", x"0F00", x"5C00", x"6B00", x"2D00", x"EFFF", x"3600", x"8100", x"4800", x"4700", x"8D00", x"9E00", x"7B00", x"AC00", x"EE00", x"A100", x"3D00", x"1200", x"D8FF", x"D5FF", x"D7FF", x"C8FF", x"9AFF", x"6BFF", x"4BFF", x"2BFF", x"34FF", x"6EFF", x"9FFF", x"B6FF", x"8EFF", x"5AFF", x"84FF", x"E3FF", x"5C00", x"A200", x"5900", x"1D00", x"0400", x"3800", x"7100", x"5A00", x"6C00", x"A000", x"A700", x"7000", x"2000", x"3E00", x"4000", x"1D00", x"0400", x"CAFF", x"C8FF", x"FBFF", x"1200", x"1200", x"C6FF", x"41FF", x"06FF", x"16FF", x"7FFF", x"C5FF", x"D0FF", x"E2FF", x"F8FF", x"DEFF", x"D7FF", x"4300", x"9600", x"B200", x"AE00", x"7600", x"4C00", x"2A00", x"1A00", x"0C00", x"1400", x"3500", x"2600", x"1C00", x"2600", x"1500", x"3900", x"5300", x"1300", x"E4FF", x"CDFF", x"E0FF", x"D6FF", x"A7FF", x"B0FF", x"7EFF", x"4BFF", x"52FF", x"74FF", x"96FF", x"C0FF", x"1D00", x"3700", x"4E00", x"5B00", x"6000", x"7A00", x"8200", x"5300", x"1700", x"2600", x"4500", x"2C00", x"1100", x"0800", x"FAFF", x"F5FF", x"0500", x"1800", x"1A00", x"1100", x"1A00", x"0700", x"D2FF", x"99FF", x"A8FF", x"BDFF", x"A6FF", x"9DFF", x"A6FF", x"A7FF", x"97FF", x"C9FF", x"FFFF", x"F6FF", x"1900", x"4200", x"4C00", x"2A00", x"1900", x"4C00", x"6A00", x"6500", x"4000", x"2D00", x"3800", x"2600", x"0B00", x"E5FF", x"B9FF", x"B1FF", x"BAFF", x"C0FF", x"D3FF", x"F0FF", x"FEFF", x"0600", x"0A00", x"FEFF", x"0200", x"1C00", x"1900", x"0900", x"F8FF", x"EFFF", x"D3FF", x"C4FF", x"D3FF", x"DDFF", x"F2FF", x"1100", x"2200", x"3100", x"5100", x"8300", x"9B00", x"7800", x"4100", x"0A00", x"E8FF", x"DDFF", x"DBFF", x"D6FF", x"B8FF", x"AEFF", x"A9FF", x"94FF", x"A9FF", x"CBFF", x"EAFF", x"FFFF", x"0000", x"2100", x"2400", x"0500", x"F3FF", x"F5FF", x"FEFF", x"F0FF", x"FBFF", x"0B00", x"1800", x"2400", x"2600", x"2A00", x"3200", x"4C00", x"6300", x"5300", x"3800", x"1500", x"0A00", x"0100", x"EBFF", x"D7FF", x"DAFF", x"D6FF", x"B9FF", x"A5FF", x"AAFF", x"B3FF", x"BAFF", x"C4FF", x"D0FF", x"DEFF", x"F5FF", x"0C00", x"1800", x"0B00", x"FDFF", x"0100", x"1600", x"2D00", x"3700", x"2E00", x"2900", x"2300", x"1200", x"0800", x"0B00", x"1100", x"1600", x"1400", x"0E00", x"0600", x"F7FF", x"F5FF", x"0000", x"FFFF", x"EFFF", x"DEFF", x"E1FF", x"EBFF", x"E1FF", x"D9FF", x"E5FF", x"F9FF", x"F7FF", x"E9FF", x"EFFF", x"0800", x"2400", x"2A00", x"3000", x"3C00", x"3700", x"1300", x"0000", x"1600", x"1D00", x"0F00", x"0900", x"0800", x"FFFF", x"FAFF", x"FDFF", x"0300", x"0400", x"0100", x"FFFF", x"0200", x"F1FF", x"D5FF", x"C2FF", x"C7FF", x"DAFF", x"E2FF", x"E0FF", x"E7FF", x"F3FF", x"F7FF", x"0100", x"1200", x"1C00", x"2200", x"2F00", x"3600", x"2000", x"0800", x"1000", x"1600", x"0500", x"F6FF", x"FAFF", x"0600", x"0100", x"F9FF", x"F1FF", x"F5FF", x"F5FF", x"F0FF", x"FCFF", x"0300", x"0500", x"0100", x"F7FF", x"F0FF", x"EAFF", x"E2FF", x"E7FF", x"F8FF", x"F8FF", x"F1FF", x"F4FF", x"0300", x"1400", x"1D00", x"1C00", x"1200", x"0F00", x"0E00", x"0700", x"FFFF", x"0300", x"0700", x"FEFF", x"F7FF", x"F5FF", x"F2FF", x"F4FF", x"EFFF", x"F7FF", x"0700", x"0B00", x"0100", x"F6FF", x"F9FF", x"FAFF", x"F9FF", x"FDFF", x"FEFF", x"0200", x"0200", x"FCFF", x"F7FF", x"F4FF", x"0100", x"1000", x"1200", x"0B00", x"0D00", x"1300", x"1400", x"0C00", x"0D00", x"1300", x"1000", x"0F00", x"0F00", x"0A00", x"0100", x"F8FF", x"F0FF", x"EFFF", x"EFFF", x"EEFF", x"F5FF", x"FDFF", x"FDFF", x"F6FF", x"F2FF", x"FAFF", x"FFFF", x"FCFF", x"FFFF", x"FFFF", x"F8FF", x"F4FF", x"F6FF", x"FAFF", x"F9FF", x"FBFF", x"FFFF", x"0500", x"0700", x"0800", x"1000", x"1700", x"1100", x"0900", x"0A00", x"0300", x"FDFF", x"0600", x"0800", x"FCFF", x"EFFF", x"F2FF", x"FCFF", x"FCFF", x"F6FF", x"F8FF", x"FBFF", x"F9FF", x"FFFF", x"0400", x"0100", x"F9FF", x"F8FF", x"FCFF", x"FFFF", x"0000", x"0500", x"0800", x"0400", x"FCFF", x"FFFF", x"0400", x"0600", x"0B00", x"1000", x"1200", x"1600", x"1100", x"0600", x"0100", x"FFFF", x"FEFF", x"FAFF", x"FAFF", x"FBFF", x"F6FF", x"EEFF", x"EBFF", x"EFFF", x"F2FF", x"F7FF", x"FEFF", x"FCFF", x"FDFF", x"0400", x"0A00", x"0800", x"0200", x"0300", x"0800", x"0600", x"FEFF", x"0000", x"0600", x"0700", x"0200", x"0400", x"0A00", x"0600", x"0000", x"FFFF", x"FFFF", x"FFFF", x"0200", x"0300", x"0100", x"FBFF", x"F7FF", x"F7FF", x"F9FF", x"F8FF", x"F7FF", x"F6FF", x"F5FF", x"F7FF", x"FEFF", x"0200", x"0200", x"0100", x"0400", x"0C00", x"0900", x"0800", x"0A00", x"0A00", x"0700", x"0300", x"0400", x"0000", x"FDFF", x"FCFF", x"FCFF", x"FCFF", x"FEFF", x"FEFF", x"FEFF", x"FFFF", x"FFFF", x"FFFF", x"FDFF", x"FCFF", x"FDFF", x"FDFF", x"FAFF", x"FEFF", x"0200", x"0000", x"0000", x"0300", x"0800", x"0200", x"FDFF", x"0000", x"0500", x"0200", x"0000", x"0100", x"0100", x"0400", x"0300", x"FFFF", x"FDFF", x"FAFF", x"FBFF", x"0000", x"0200", x"0300", x"0100", x"0400", x"0400", x"0100", x"0000", x"FEFF", x"0000", x"FEFF", x"FDFF", x"0000", x"0200", x"0300", x"0600", x"0700", x"0600", x"0500", x"0600", x"0200", x"0400", x"0400", x"0000", x"0100", x"FFFF", x"FDFF", x"FBFF", x"FDFF", x"0100", x"0100", x"0000", x"FFFF", x"0000", x"FCFF", x"FBFF", x"0000", x"0000", x"FDFF", x"FDFF", x"FEFF", x"FEFF", x"FBFF", x"FDFF", x"0100", x"0300", x"0000", x"FFFF", x"0300", x"0100", x"FEFF", x"FBFF", x"FDFF", x"FCFF", x"FBFF", x"FEFF", x"0100", x"FFFF", x"FDFF", x"FFFF", x"FFFF", x"FFFF", x"0000", x"0000", x"FEFF", x"FEFF", x"0100", x"0100", x"FFFF", x"0000", x"FFFF", x"FCFF", x"FBFF", x"FBFF", x"FEFF", x"FEFF", x"0100", x"0300", x"0400", x"0400", x"0400", x"0400", x"0100", x"0200", x"0300", x"0200", x"FFFF", x"0000", x"0400", x"0200", x"0300", x"0400", x"0300", x"0000", x"FBFF", x"FCFF", x"FCFF", x"FEFF", x"FDFF", x"FCFF", x"FCFF", x"FDFF", x"FDFF", x"0000", x"0200", x"0200", x"0300", x"0300", x"0400", x"0200", x"0300", x"0400", x"0400", x"0500", x"0400", x"0300", x"0400", x"0200", x"0100", x"0200", x"0200", x"0300", x"0500", x"0400", x"0100", x"0100", x"0000", x"0200", x"FEFF", x"FFFF", x"FFFF", x"FDFF", x"FEFF", x"FDFF", x"FDFF", x"FBFF", x"F9FF", x"FCFF", x"0000", x"0100", x"FFFF", x"0000", x"0200", x"FFFF", x"FFFF", x"0100", x"0100", x"0000", x"0000", x"0300", x"0300", x"0000", x"0100", x"FEFF", x"FDFF", x"FDFF", x"FBFF", x"F9FF", x"FCFF", x"FEFF", x"0100", x"FFFF", x"FEFF", x"0000", x"0000", x"0000", x"FFFF", x"FCFF", x"F9FF", x"F9FF", x"F9FF", x"F8FF", x"FCFF", x"FCFF", x"FCFF", x"FEFF", x"0100", x"0200", x"0200", x"0400", x"0300", x"0200", x"0400", x"0300", x"0500", x"0600", x"0800", x"0700", x"0500", x"0600", x"0500", x"0300", x"0400", x"0400", x"0300", x"0400", x"0300", x"0100", x"0300", x"0100", x"0000", x"0200", x"0300", x"0000", x"FEFF", x"FFFF", x"FEFF", x"FFFF", x"FDFF", x"FDFF", x"FDFF", x"FDFF", x"FEFF", x"FFFF", x"FFFF", x"FDFF", x"FEFF", x"0000", x"FFFF", x"FEFF", x"0000", x"0000", x"0200", x"0400", x"0200", x"0300", x"0200", x"0000", x"FFFF", x"FFFF", x"FFFF", x"FBFF", x"FCFF", x"FAFF", x"FAFF", x"FCFF", x"FDFF", x"FFFF", x"0100", x"0100", x"0100", x"0200", x"0300", x"0200", x"0300", x"0400", x"0400", x"0300", x"0400", x"FFFF", x"FCFF", x"FBFF", x"FCFF", x"FFFF", x"FFFF", x"0000", x"FFFF", x"0100", x"0100", x"0100", x"0200", x"0200", x"0200", x"0100", x"0000", x"FFFF", x"FEFF", x"FEFF", x"FEFF", x"FEFF", x"FEFF", x"FDFF", x"FCFF", x"FDFF", x"FFFF", x"FEFF", x"0000", x"FFFF", x"FEFF", x"FDFF", x"FDFF", x"FDFF", x"FCFF", x"FEFF", x"0100", x"0100", x"0100", x"0200", x"0200", x"0100", x"0300", x"0300", x"FFFF", x"0100", x"0200", x"0300", x"0500", x"0200", x"0200", x"0200", x"0200", x"0300", x"0100", x"0200", x"0300", x"0200", x"0200", x"0000", x"FFFF", x"FFFF", x"FFFF", x"0100", x"0100", x"0200", x"0100", x"0000", x"0000", x"0100", x"0100", x"0100", x"0300", x"0200", x"FFFF", x"0000", x"FDFF", x"FAFF", x"FEFF", x"FFFF", x"FDFF", x"FDFF", x"FEFF", x"FFFF", x"FDFF", x"FCFF", x"FDFF", x"FEFF", x"FFFF", x"0100", x"0200", x"0400", x"0200", x"0300", x"0300", x"0400", x"0600", x"0300", x"0200", x"0100", x"0200", x"0200", x"0000", x"0100", x"FFFF", x"0000", x"0100", x"0000", x"0200", x"0200", x"FFFF", x"FEFF", x"FEFF", x"FBFF", x"FDFF", x"FDFF", x"FDFF", x"FEFF", x"FEFF", x"FDFF", x"FDFF", x"FFFF", x"0100", x"0100", x"0000", x"FFFF", x"FCFF", x"FDFF", x"0000", x"FFFF", x"FDFF", x"FBFF", x"FDFF", x"FEFF", x"FDFF", x"FEFF", x"FEFF", x"FEFF", x"0000", x"0200", x"0300", x"0200", x"0100", x"0000", x"0000", x"FEFF", x"0200", x"0200", x"0200", x"0000", x"0000", x"0100", x"0000", x"0200", x"0200", x"0100", x"FFFF", x"FCFF", x"FEFF", x"FEFF", x"0000", x"0000", x"0200", x"0400", x"0300", x"0200", x"FEFF", x"0200", x"0300", x"0200", x"0200", x"0200", x"0400", x"0400", x"0300", x"0300", x"0300", x"0500", x"0600", x"0500", x"0500", x"0300", x"0400", x"0100", x"0100", x"0100", x"0100", x"0100", x"FFFF", x"FFFF", x"0000", x"FFFF", x"FEFF", x"FCFF", x"0000", x"FFFF", x"FEFF", x"0000", x"FFFF", x"FFFF", x"FEFF", x"FEFF", x"FDFF", x"FDFF", x"FCFF", x"F9FF", x"FAFF", x"FBFF", x"FBFF", x"FDFF", x"FCFF", x"FAFF", x"FCFF", x"FCFF", x"FAFF", x"FBFF", x"FBFF", x"FDFF", x"FEFF", x"0200", x"0000", x"0000", x"0000", x"FCFF", x"0000", x"0100", x"0200", x"0200", x"0000", x"0100", x"0100", x"0400", x"0400", x"0300", x"0300", x"0400", x"0600", x"0400", x"0300", x"0200", x"0400", x"0300", x"0200", x"0200", x"0200", x"0100", x"0000", x"0200", x"0400", x"0400", x"0300", x"0300", x"0200", x"0100", x"0000", x"0300", x"0000", x"0000", x"FFFF", x"FEFF", x"0000", x"FEFF", x"0100", x"FEFF", x"FCFF", x"FFFF", x"FDFF", x"FEFF", x"0000", x"0000", x"0100", x"FFFF", x"0300", x"0100", x"FFFF", x"0000", x"FDFF", x"FDFF", x"FDFF", x"FFFF", x"FFFF", x"FDFF", x"FFFF", x"FEFF", x"FDFF", x"FEFF", x"FCFF", x"FCFF", x"FCFF", x"FDFF", x"FEFF", x"0000", x"0200", x"0200", x"0200", x"0400", x"0100", x"0000", x"FFFF", x"FFFF", x"FDFF", x"FEFF", x"0000", x"0100", x"0100", x"0100", x"0100", x"0100", x"0200", x"0200", x"0100", x"FDFF", x"FEFF", x"0000", x"0000", x"0100", x"0100", x"FFFF", x"0000", x"0100", x"0200", x"0400", x"0300", x"0400", x"0400", x"0500", x"0400", x"0400", x"0200", x"0000", x"0100", x"0100", x"0300", x"0300", x"0400", x"0200", x"0200", x"0200", x"0100", x"0100", x"0200", x"0300", x"0000", x"FFFF", x"FEFF", x"FEFF", x"FEFF", x"FDFF", x"FDFF", x"FDFF", x"FDFF", x"0000", x"0100", x"0200", x"0000", x"FEFF", x"0100", x"FFFF", x"0000", x"FEFF", x"FEFF", x"FFFF", x"FDFF", x"FCFF", x"FAFF", x"FBFF", x"FDFF", x"FDFF", x"FFFF", x"FFFF", x"0300", x"FEFF", x"0600", x"0400", x"F9FF", x"EBFF", x"F4FF", x"0000", x"FAFF", x"0400", x"0500");
				--
				signal Bes_voice : Bes :=(x"494E", x"464F", x"4953", x"4654", x"0E00", x"0000", x"4C61", x"7666", x"3538", x"2E37", x"362E", x"3130", x"3000", x"6461", x"7461", x"4824", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"FFFF", x"0000", x"0100", x"0000", x"0000", x"0000", x"0100", x"0000", x"0000", x"0000", x"FFFF", x"0100", x"0000", x"FFFF", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"FFFF", x"FEFF", x"0100", x"0000", x"FCFF", x"FEFF", x"0000", x"FEFF", x"0200", x"0000", x"0400", x"0600", x"0500", x"0300", x"FEFF", x"0300", x"0600", x"0200", x"0500", x"0600", x"0100", x"0000", x"FEFF", x"FEFF", x"FFFF", x"FDFF", x"0000", x"0400", x"0200", x"0500", x"0500", x"0600", x"0200", x"FDFF", x"FFFF", x"FBFF", x"F8FF", x"F4FF", x"F5FF", x"F6FF", x"FBFF", x"FDFF", x"FBFF", x"0300", x"0600", x"0500", x"0600", x"0900", x"0800", x"0400", x"0400", x"0200", x"FCFF", x"F9FF", x"FEFF", x"0000", x"0300", x"0600", x"0200", x"0100", x"0400", x"0600", x"0400", x"0400", x"0500", x"0400", x"0200", x"0100", x"FEFF", x"FCFF", x"FCFF", x"FDFF", x"FCFF", x"FDFF", x"FFFF", x"FFFF", x"FEFF", x"FEFF", x"0100", x"0100", x"FEFF", x"FDFF", x"FEFF", x"FBFF", x"FBFF", x"FDFF", x"FBFF", x"FAFF", x"FDFF", x"FDFF", x"FAFF", x"FCFF", x"FCFF", x"FCFF", x"0500", x"0700", x"0700", x"0900", x"0A00", x"0A00", x"0200", x"0100", x"0100", x"0000", x"FBFF", x"F8FF", x"FDFF", x"FDFF", x"FBFF", x"FFFF", x"FFFF", x"FDFF", x"FDFF", x"FFFF", x"0400", x"FEFF", x"FEFF", x"FFFF", x"0000", x"0000", x"FFFF", x"0300", x"0000", x"0000", x"0100", x"0100", x"FCFF", x"FEFF", x"0100", x"0000", x"0000", x"0200", x"0100", x"FFFF", x"0200", x"0300", x"0200", x"0300", x"0600", x"0900", x"0800", x"0900", x"0900", x"0700", x"0300", x"0100", x"0000", x"FFFF", x"FEFF", x"FCFF", x"FBFF", x"FCFF", x"FDFF", x"FEFF", x"0100", x"0200", x"0300", x"0500", x"0400", x"0100", x"FFFF", x"FDFF", x"FDFF", x"FAFF", x"FBFF", x"F9FF", x"F8FF", x"F6FF", x"F6FF", x"FAFF", x"FDFF", x"FCFF", x"FDFF", x"FDFF", x"FFFF", x"0000", x"0000", x"FFFF", x"FCFF", x"0100", x"0300", x"0300", x"FDFF", x"0200", x"0400", x"0300", x"0B00", x"0C00", x"0B00", x"0700", x"0400", x"0200", x"0300", x"0100", x"0200", x"0000", x"FCFF", x"F8FF", x"FEFF", x"FDFF", x"FEFF", x"0200", x"0100", x"0000", x"FFFF", x"FDFF", x"FEFF", x"0100", x"0100", x"0100", x"FEFF", x"FAFF", x"FBFF", x"FAFF", x"FCFF", x"0100", x"0000", x"0300", x"0200", x"0400", x"0600", x"0500", x"0300", x"0200", x"0400", x"0300", x"0100", x"0200", x"0200", x"FFFF", x"0100", x"0000", x"FCFF", x"F8FF", x"F7FF", x"F8FF", x"FCFF", x"F9FF", x"FFFF", x"0100", x"FFFF", x"FFFF", x"0000", x"0400", x"0300", x"FFFF", x"FFFF", x"0100", x"0200", x"FFFF", x"0400", x"0400", x"0300", x"0500", x"0400", x"0100", x"FDFF", x"FFFF", x"FDFF", x"F9FF", x"FBFF", x"F9FF", x"FCFF", x"FFFF", x"0300", x"0500", x"0100", x"FFFF", x"0100", x"0200", x"0100", x"0100", x"0100", x"FEFF", x"FAFF", x"0000", x"0100", x"0400", x"0300", x"0600", x"0300", x"FFFF", x"0200", x"0200", x"0100", x"0300", x"0500", x"0700", x"0700", x"0100", x"0400", x"0100", x"FBFF", x"FBFF", x"F8FF", x"F9FF", x"F6FF", x"F9FF", x"FCFF", x"FCFF", x"FBFF", x"FDFF", x"0200", x"0000", x"FAFF", x"FBFF", x"FDFF", x"0000", x"0400", x"0300", x"0800", x"0400", x"0400", x"0500", x"0200", x"FFFF", x"0000", x"FFFF", x"0200", x"0000", x"0200", x"0400", x"0100", x"0200", x"0300", x"0700", x"0300", x"0300", x"0100", x"FFFF", x"FDFF", x"FAFF", x"F9FF", x"FDFF", x"FBFF", x"FEFF", x"0500", x"0300", x"0300", x"0200", x"0000", x"0200", x"0000", x"FEFF", x"FDFF", x"FBFF", x"FFFF", x"0000", x"FCFF", x"FBFF", x"FFFF", x"FEFF", x"FEFF", x"FDFF", x"FDFF", x"FDFF", x"FDFF", x"FDFF", x"FBFF", x"FBFF", x"FCFF", x"F8FF", x"FAFF", x"FCFF", x"FEFF", x"0000", x"FFFF", x"FFFF", x"0200", x"0100", x"FFFF", x"0700", x"0900", x"0500", x"0A00", x"0F00", x"0800", x"0800", x"0A00", x"0B00", x"0900", x"0200", x"0600", x"0600", x"0600", x"0800", x"0400", x"0100", x"0300", x"0200", x"0000", x"FCFF", x"0000", x"0000", x"FAFF", x"FDFF", x"FBFF", x"F8FF", x"FAFF", x"FBFF", x"FBFF", x"FBFF", x"FAFF", x"FCFF", x"FEFF", x"FEFF", x"0100", x"FFFF", x"0000", x"0600", x"0300", x"0500", x"0500", x"0200", x"0000", x"FEFF", x"0000", x"FDFF", x"FBFF", x"FDFF", x"F9FF", x"F7FF", x"FBFF", x"FEFF", x"0000", x"0300", x"0400", x"0400", x"0300", x"0500", x"0400", x"0200", x"FFFF", x"F9FF", x"FAFF", x"FAFF", x"F8FF", x"FEFF", x"0300", x"0000", x"0000", x"0200", x"FAFF", x"FCFF", x"FFFF", x"FBFF", x"F8FF", x"FAFF", x"FDFF", x"FEFF", x"0100", x"0500", x"0400", x"FCFF", x"FBFF", x"FBFF", x"FAFF", x"FDFF", x"FFFF", x"0000", x"0200", x"0300", x"0400", x"0600", x"0A00", x"0B00", x"0D00", x"0D00", x"0A00", x"0B00", x"0900", x"0A00", x"0600", x"0400", x"0300", x"FEFF", x"0100", x"FDFF", x"FAFF", x"FAFF", x"FFFF", x"0000", x"0200", x"0600", x"0500", x"0100", x"0100", x"FDFF", x"FAFF", x"FBFF", x"FEFF", x"FDFF", x"FAFF", x"FBFF", x"FCFF", x"FDFF", x"FCFF", x"FCFF", x"FFFF", x"0000", x"0400", x"0300", x"0100", x"FFFF", x"FAFF", x"F9FF", x"F6FF", x"F6FF", x"FCFF", x"FDFF", x"0000", x"FFFF", x"FCFF", x"FCFF", x"FFFF", x"F9FF", x"F9FF", x"FCFF", x"FEFF", x"0000", x"FFFF", x"FEFF", x"FFFF", x"0100", x"0300", x"0200", x"0000", x"0300", x"0700", x"0700", x"0700", x"0700", x"0600", x"0300", x"0400", x"0300", x"0500", x"0600", x"0200", x"0400", x"0400", x"0400", x"0700", x"0700", x"0600", x"0300", x"0300", x"0100", x"FCFF", x"FAFF", x"FEFF", x"FFFF", x"FFFF", x"0400", x"0300", x"0200", x"0300", x"0100", x"FDFF", x"FBFF", x"FCFF", x"FEFF", x"0100", x"FBFF", x"FCFF", x"FCFF", x"0000", x"0300", x"0200", x"FFFF", x"FEFF", x"0300", x"0100", x"0200", x"0100", x"0300", x"0300", x"FCFF", x"FDFF", x"FEFF", x"FBFF", x"F6FF", x"FAFF", x"FCFF", x"FDFF", x"FFFF", x"FFFF", x"FDFF", x"FDFF", x"0000", x"FCFF", x"FDFF", x"FBFF", x"F8FF", x"F9FF", x"F9FF", x"F8FF", x"F9FF", x"FAFF", x"FDFF", x"0000", x"FFFF", x"0200", x"0500", x"0400", x"0300", x"0500", x"0500", x"0400", x"0000", x"0100", x"0300", x"0800", x"0C00", x"0C00", x"1000", x"0A00", x"0600", x"0500", x"0600", x"0800", x"0300", x"0200", x"0300", x"0500", x"0300", x"0200", x"0300", x"FBFF", x"F9FF", x"FAFF", x"FAFF", x"FCFF", x"FDFF", x"FBFF", x"FDFF", x"FEFF", x"FCFF", x"FBFF", x"FAFF", x"FDFF", x"FEFF", x"FFFF", x"FFFF", x"FDFF", x"FFFF", x"FCFF", x"FFFF", x"FEFF", x"FFFF", x"FDFF", x"FBFF", x"FEFF", x"FCFF", x"0300", x"0400", x"0500", x"0500", x"0600", x"0400", x"0400", x"0400", x"0200", x"0100", x"0000", x"FFFF", x"FBFF", x"0000", x"0200", x"FDFF", x"0200", x"0200", x"FFFF", x"FDFF", x"FBFF", x"0200", x"0500", x"0400", x"0000", x"FFFF", x"FDFF", x"FCFF", x"FCFF", x"FAFF", x"FBFF", x"F7FF", x"FAFF", x"0100", x"0400", x"0800", x"0700", x"FFFF", x"0100", x"0300", x"FFFF", x"FEFF", x"FEFF", x"0100", x"0300", x"0500", x"0300", x"0200", x"FCFF", x"FAFF", x"F6FF", x"F7FF", x"F6FF", x"F7FF", x"0100", x"0400", x"0500", x"0500", x"0100", x"0000", x"FDFF", x"FEFF", x"FFFF", x"FEFF", x"FAFF", x"FBFF", x"FEFF", x"FEFF", x"FFFF", x"0300", x"0700", x"0400", x"0700", x"0600", x"0400", x"0500", x"0000", x"0300", x"0200", x"0700", x"0400", x"0500", x"0400", x"0300", x"0400", x"0400", x"FEFF", x"0200", x"0300", x"0400", x"0800", x"0400", x"0100", x"FEFF", x"FFFF", x"FDFF", x"FEFF", x"0200", x"0100", x"0300", x"0300", x"0000", x"FDFF", x"FEFF", x"FEFF", x"FAFF", x"FAFF", x"FAFF", x"FAFF", x"FEFF", x"0200", x"0200", x"0100", x"0000", x"0200", x"0000", x"FCFF", x"FEFF", x"FCFF", x"F9FF", x"F6FF", x"F9FF", x"F8FF", x"FCFF", x"FEFF", x"0200", x"0300", x"0100", x"0100", x"0600", x"0400", x"0200", x"0400", x"0100", x"0200", x"0200", x"0200", x"0700", x"0800", x"0800", x"0300", x"0100", x"0100", x"0300", x"0300", x"FEFF", x"0100", x"0200", x"FEFF", x"0100", x"FFFF", x"FCFF", x"F5FF", x"F5FF", x"F6FF", x"F6FF", x"F9FF", x"F8FF", x"FBFF", x"FCFF", x"FFFF", x"FDFF", x"FFFF", x"FEFF", x"0000", x"0100", x"0300", x"0100", x"FCFF", x"FFFF", x"FDFF", x"FEFF", x"FCFF", x"FBFF", x"FDFF", x"0200", x"0600", x"0500", x"0800", x"0800", x"0600", x"0300", x"0400", x"FEFF", x"0200", x"0600", x"0600", x"0400", x"0200", x"0400", x"0400", x"0300", x"0000", x"0000", x"FDFF", x"0000", x"0500", x"0300", x"0600", x"FFFF", x"FCFF", x"FBFF", x"FAFF", x"FBFF", x"FEFF", x"FFFF", x"0100", x"0200", x"FDFF", x"FFFF", x"0000", x"FCFF", x"0000", x"0000", x"FEFF", x"FFFF", x"FEFF", x"FEFF", x"FAFF", x"FDFF", x"FDFF", x"0100", x"0400", x"0400", x"0600", x"0200", x"0100", x"0100", x"FFFF", x"FBFF", x"FCFF", x"0100", x"0200", x"0200", x"0000", x"0500", x"0500", x"0300", x"0300", x"0200", x"0700", x"0500", x"0300", x"FFFF", x"FCFF", x"FBFF", x"FBFF", x"FCFF", x"0200", x"FCFF", x"FAFF", x"FAFF", x"F9FF", x"FCFF", x"FEFF", x"FDFF", x"FEFF", x"0500", x"0400", x"0300", x"0900", x"0B00", x"0700", x"0400", x"0400", x"0300", x"0500", x"0700", x"0800", x"0900", x"0600", x"0600", x"0900", x"0700", x"0600", x"0700", x"0200", x"FEFF", x"FBFF", x"FBFF", x"F9FF", x"F8FF", x"F6FF", x"F7FF", x"F8FF", x"FAFF", x"FDFF", x"FDFF", x"FFFF", x"FFFF", x"FFFF", x"0200", x"0100", x"0100", x"0200", x"0600", x"0200", x"FEFF", x"FBFF", x"F5FF", x"F5FF", x"F7FF", x"F8FF", x"F7FF", x"F7FF", x"F2FF", x"F3FF", x"F7FF", x"F9FF", x"FDFF", x"FBFF", x"0300", x"0200", x"0100", x"0400", x"0300", x"0400", x"0600", x"0700", x"0500", x"0700", x"0600", x"0000", x"0700", x"0800", x"0800", x"0800", x"0800", x"0300", x"0000", x"FDFF", x"F8FF", x"F9FF", x"0000", x"0200", x"0400", x"0600", x"0700", x"0300", x"0200", x"0300", x"FFFF", x"FFFF", x"FEFF", x"F9FF", x"FBFF", x"FAFF", x"FDFF", x"0000", x"0100", x"0200", x"0500", x"0600", x"0700", x"0800", x"0600", x"0200", x"0100", x"FEFF", x"F7FF", x"F8FF", x"F7FF", x"F9FF", x"F9FF", x"FBFF", x"0000", x"0000", x"FFFF", x"FEFF", x"FDFF", x"FEFF", x"FCFF", x"F9FF", x"F5FF", x"F9FF", x"FEFF", x"FEFF", x"0300", x"0700", x"0900", x"0500", x"0A00", x"0B00", x"0700", x"0900", x"0300", x"0000", x"0200", x"0200", x"0300", x"0600", x"0500", x"0600", x"0500", x"0100", x"0400", x"FFFF", x"0000", x"0100", x"0100", x"0100", x"FEFF", x"FFFF", x"FDFF", x"FEFF", x"FDFF", x"FDFF", x"FEFF", x"FDFF", x"FBFF", x"F9FF", x"FAFF", x"FBFF", x"FEFF", x"0000", x"0000", x"0200", x"0300", x"0100", x"0100", x"FFFF", x"0100", x"FFFF", x"0100", x"0100", x"FEFF", x"0200", x"FCFF", x"FCFF", x"FDFF", x"0000", x"0200", x"0400", x"0700", x"0800", x"0300", x"FFFF", x"FDFF", x"FBFF", x"F7FF", x"F7FF", x"FAFF", x"F9FF", x"FBFF", x"FDFF", x"0000", x"FFFF", x"0000", x"0100", x"0000", x"FFFF", x"0000", x"FEFF", x"FFFF", x"FCFF", x"FBFF", x"F9FF", x"F8FF", x"FBFF", x"F9FF", x"F9FF", x"FBFF", x"FAFF", x"FDFF", x"0100", x"0400", x"0700", x"0700", x"0900", x"0D00", x"0D00", x"0D00", x"0700", x"0500", x"0500", x"0100", x"0200", x"FFFF", x"FDFF", x"FCFF", x"FDFF", x"0200", x"0300", x"0800", x"0A00", x"0800", x"0600", x"0400", x"0100", x"FFFF", x"FFFF", x"FEFF", x"0300", x"0600", x"0600", x"0400", x"0100", x"0400", x"0800", x"0400", x"0800", x"0300", x"FEFF", x"0100", x"0100", x"0000", x"0300", x"FEFF", x"0100", x"0000", x"FBFF", x"FCFF", x"FBFF", x"FEFF", x"FEFF", x"F9FF", x"FBFF", x"FCFF", x"F7FF", x"F6FF", x"FBFF", x"FAFF", x"F8FF", x"F9FF", x"F9FF", x"F8FF", x"F6FF", x"FDFF", x"FCFF", x"FDFF", x"FDFF", x"0200", x"0000", x"0000", x"0100", x"FEFF", x"FFFF", x"0000", x"FFFF", x"FEFF", x"0100", x"0300", x"0300", x"0600", x"0800", x"0600", x"0800", x"0400", x"0200", x"0600", x"0700", x"0B00", x"0900", x"0800", x"0400", x"FDFF", x"FBFF", x"FBFF", x"FAFF", x"FDFF", x"FDFF", x"FBFF", x"F8FF", x"FBFF", x"FBFF", x"F7FF", x"FCFF", x"FAFF", x"FCFF", x"FEFF", x"0000", x"FFFF", x"FFFF", x"0200", x"0000", x"FBFF", x"FAFF", x"FBFF", x"FEFF", x"0300", x"0500", x"0700", x"0800", x"0800", x"0800", x"0900", x"0900", x"0900", x"0700", x"0600", x"0200", x"0000", x"FEFF", x"FDFF", x"FDFF", x"FCFF", x"FDFF", x"0000", x"FFFF", x"0100", x"FEFF", x"FFFF", x"0300", x"0000", x"FEFF", x"FEFF", x"FDFF", x"FBFF", x"FAFF", x"F7FF", x"FEFF", x"0200", x"0500", x"0700", x"0300", x"0300", x"0500", x"0800", x"0200", x"0000", x"0200", x"FCFF", x"FBFF", x"FCFF", x"FEFF", x"FEFF", x"0000", x"0300", x"0100", x"0000", x"0000", x"0000", x"0000", x"FFFF", x"0300", x"0500", x"0500", x"0600", x"0700", x"0400", x"0300", x"FFFF", x"FAFF", x"FEFF", x"FEFF", x"0000", x"FDFF", x"FEFF", x"FFFF", x"FDFF", x"FEFF", x"FAFF", x"F8FF", x"FAFF", x"FDFF", x"FDFF", x"FDFF", x"0000", x"0200", x"0100", x"0400", x"0200", x"0100", x"FFFF", x"0300", x"0400", x"0100", x"0500", x"0900", x"0800", x"0900", x"0900", x"0300", x"FFFF", x"FFFF", x"FCFF", x"F9FF", x"F9FF", x"F5FF", x"F4FF", x"F4FF", x"F7FF", x"F8FF", x"FAFF", x"FAFF", x"0100", x"0400", x"0700", x"0300", x"0100", x"0200", x"0100", x"FEFF", x"FDFF", x"FBFF", x"FDFF", x"FDFF", x"FFFF", x"0000", x"0200", x"0300", x"0200", x"0600", x"0300", x"0400", x"0500", x"0600", x"0000", x"0000", x"FEFF", x"FAFF", x"0100", x"0100", x"FCFF", x"0200", x"0200", x"0000", x"0100", x"0300", x"0200", x"0500", x"0700", x"0A00", x"0700", x"0400", x"0100", x"0000", x"0100", x"0000", x"FDFF", x"0000", x"0100", x"FFFF", x"FFFF", x"FFFF", x"0100", x"FEFF", x"0000", x"0000", x"0100", x"0200", x"0000", x"0100", x"0100", x"0000", x"FBFF", x"FBFF", x"FAFF", x"FBFF", x"FAFF", x"FFFF", x"0200", x"0200", x"0100", x"FEFF", x"FCFF", x"FCFF", x"FDFF", x"FBFF", x"FDFF", x"FEFF", x"0000", x"0500", x"0700", x"0400", x"0600", x"0400", x"FDFF", x"0000", x"FFFF", x"FCFF", x"FDFF", x"FEFF", x"FEFF", x"0200", x"0400", x"0400", x"FFFF", x"0200", x"0000", x"FDFF", x"FDFF", x"F9FF", x"FEFF", x"FDFF", x"FDFF", x"FFFF", x"0000", x"FFFF", x"FEFF", x"FEFF", x"0300", x"0300", x"0300", x"0000", x"FFFF", x"FDFF", x"FFFF", x"0100", x"FEFF", x"0100", x"0400", x"0800", x"0400", x"0100", x"FEFF", x"0100", x"0000", x"FDFF", x"0100", x"0200", x"0000", x"0000", x"0100", x"0200", x"0000", x"FEFF", x"0000", x"0100", x"0500", x"0B00", x"0D00", x"0A00", x"0600", x"0100", x"FEFF", x"FFFF", x"FFFF", x"FDFF", x"FFFF", x"FFFF", x"FFFF", x"0500", x"0100", x"FDFF", x"F7FF", x"F5FF", x"F6FF", x"F7FF", x"F8FF", x"FDFF", x"FDFF", x"0200", x"0500", x"0200", x"0300", x"0200", x"0500", x"0400", x"0400", x"0100", x"FFFF", x"0000", x"FFFF", x"0000", x"FEFF", x"FBFF", x"F9FF", x"FDFF", x"FFFF", x"FBFF", x"FEFF", x"FCFF", x"FFFF", x"0600", x"0100", x"0100", x"0000", x"0100", x"0100", x"0300", x"0400", x"0300", x"FFFF", x"FFFF", x"0100", x"FEFF", x"0100", x"0200", x"0500", x"0600", x"0400", x"0200", x"0300", x"0300", x"FFFF", x"0100", x"FEFF", x"FFFF", x"FBFF", x"FEFF", x"0000", x"FBFF", x"FAFF", x"FAFF", x"F6FF", x"FBFF", x"FEFF", x"FCFF", x"0100", x"0100", x"FDFF", x"FEFF", x"FFFF", x"FDFF", x"FCFF", x"FFFF", x"0300", x"0100", x"0200", x"0500", x"0300", x"0700", x"0900", x"0300", x"0100", x"0000", x"FDFF", x"FBFF", x"F8FF", x"F8FF", x"FDFF", x"FDFF", x"0100", x"0500", x"0500", x"0600", x"0800", x"0900", x"0900", x"0B00", x"0C00", x"0A00", x"0900", x"0700", x"0A00", x"0B00", x"0500", x"0700", x"0200", x"FEFF", x"FBFF", x"F7FF", x"F9FF", x"F4FF", x"F5FF", x"F8FF", x"F8FF", x"F7FF", x"F9FF", x"F3FF", x"F5FF", x"F6FF", x"FBFF", x"0200", x"0800", x"0E00", x"1100", x"1300", x"1300", x"1300", x"1000", x"0700", x"0100", x"FDFF", x"F1FF", x"ECFF", x"E7FF", x"E7FF", x"E3FF", x"DEFF", x"DEFF", x"E0FF", x"E8FF", x"EFFF", x"F7FF", x"FCFF", x"0300", x"0D00", x"1300", x"1A00", x"2400", x"2800", x"2A00", x"3100", x"3600", x"3500", x"2F00", x"2700", x"2300", x"1100", x"FCFF", x"E2FF", x"C7FF", x"A9FF", x"8EFF", x"7AFF", x"73FF", x"74FF", x"84FF", x"9DFF", x"BCFF", x"E2FF", x"0B00", x"3500", x"5F00", x"8700", x"A900", x"C800", x"E200", x"F700", x"0401", x"0101", x"E900", x"AF00", x"5600", x"DFFF", x"4CFF", x"B4FE", x"1EFE", x"A2FD", x"52FD", x"39FD", x"62FD", x"CDFD", x"6AFE", x"3FFF", x"3500", x"3701", x"3602", x"0B03", x"A903", x"FD03", x"0804", x"D503", x"5B03", x"B302", x"D501", x"D200", x"BEFF", x"A6FE", x"A5FD", x"BDFC", x"FDFB", x"6BFB", x"01FB", x"CCFA", x"D1FA", x"16FB", x"A5FB", x"90FC", x"E2FD", x"86FF", x"6B01", x"4503", x"EB04", x"3206", x"E806", x"1C07", x"C406", x"EB05", x"AB04", x"0D03", x"4901", x"73FF", x"C7FD", x"81FC", x"A3FB", x"6BFB", x"BBFB", x"84FC", x"A6FD", x"D7FE", x"ECFF", x"A100", x"BE00", x"4800", x"4CFF", x"02FE", x"B9FC", x"D0FB", x"82FB", x"01FC", x"51FD", x"04FF", x"0001", x"CC02", x"4804", x"7B05", x"2806", x"7106", x"2A06", x"5205", x"1D04", x"8302", x"EA00", x"7AFF", x"53FE", x"ACFD", x"64FD", x"6FFD", x"A9FD", x"D4FD", x"DDFD", x"7CFD", x"C1FC", x"CFFB", x"D5FA", x"74FA", x"B3FA", x"E5FB", x"E7FD", x"0F00", x"6202", x"3204", x"8305", x"8006", x"DC06", x"F406", x"7506", x"7205", x"1404", x"4002", x"8200", x"E6FE", x"B8FD", x"2EFD", x"04FD", x"64FD", x"F4FD", x"7EFE", x"D9FE", x"9AFE", x"D2FD", x"7CFC", x"EFFA", x"9DF9", x"10F9", x"75F9", x"FFFA", x"59FD", x"E9FF", x"8202", x"8D04", x"2106", x"3707", x"B907", x"E107", x"5F07", x"4406", x"9604", x"5402", x"0200", x"D9FD", x"52FC", x"A7FB", x"AEFB", x"61FC", x"55FD", x"46FE", x"F1FE", x"01FF", x"70FE", x"4EFD", x"E6FB", x"BCFA", x"4BFA", x"BFFA", x"5EFC", x"7FFE", x"D900", x"0E03", x"9504", x"E705", x"B206", x"2007", x"5307", x"C306", x"CF05", x"1B04", x"0502", x"FAFF", x"11FE", x"DFFC", x"40FC", x"46FC", x"D2FC", x"72FD", x"24FE", x"71FE", x"4BFE", x"A4FD", x"8BFC", x"57FB", x"70FA", x"54FA", x"05FB", x"E4FC", x"25FF", x"8701", x"B603", x"3C05", x"8B06", x"4007", x"A507", x"AA07", x"E506", x"A205", x"A103", x"4601", x"1AFF", x"2DFD", x"0AFC", x"9AFB", x"C9FB", x"93FC", x"7EFD", x"66FE", x"E5FE", x"CCFE", x"11FE", x"CCFC", x"57FB", x"56FA", x"11FA", x"BFFA", x"B4FC", x"DDFE", x"5A01", x"8D03", x"2005", x"9506", x"6207", x"0808", x"2308", x"6007", x"1506", x"E103", x"6E01", x"20FF", x"1CFD", x"F6FB", x"5AFB", x"7FFB", x"13FC", x"C2FC", x"92FD", x"EFFD", x"EBFD", x"4EFD", x"48FC", x"23FB", x"55FA", x"56FA", x"33FB", x"3DFD", x"A8FF", x"3002", x"7E04", x"1E06", x"7D07", x"3C08", x"A408", x"8F08", x"9807", x"2406", x"D503", x"3C01", x"D2FE", x"ACFC", x"73FB", x"F8FA", x"2BFB", x"E7FB", x"BEFC", x"92FD", x"FAFD", x"EBFD", x"49FD", x"2DFC", x"D3FA", x"BEF9", x"6EF9", x"EEF9", x"D0FB", x"53FE", x"0B01", x"D903", x"DF05", x"9A07", x"C208", x"5A09", x"9D09", x"E608", x"8A07", x"7005", x"C602", x"3400", x"C6FD", x"28FC", x"3DFB", x"ECFA", x"43FB", x"A6FB", x"50FC", x"B0FC", x"BDFC", x"73FC", x"A2FB", x"C8FA", x"ECF9", x"C4F9", x"57FA", x"F1FB", x"7EFE", x"2601", x"F703", x"3B06", x"E607", x"2509", x"A509", x"C909", x"2F09", x"CC07", x"E005", x"2F03", x"7B00", x"E9FD", x"D0FB", x"9CFA", x"05FA", x"52FA", x"1AFB", x"1CFC", x"34FD", x"D2FD", x"08FE", x"A1FD", x"AAFC", x"8AFB", x"59FA", x"C3F9", x"EFF9", x"14FB", x"78FD", x"3D00", x"5803", x"2106", x"2608", x"BC09", x"790A", x"9D0A", x"1C0A", x"AF08", x"A506", x"F703", x"0F01", x"4DFE", x"F9FB", x"76FA", x"A1F9", x"A5F9", x"34FA", x"16FB", x"2FFC", x"EAFC", x"52FD", x"1DFD", x"59FC", x"51FB", x"20FA", x"5FF9", x"71F9", x"6EFA", x"A1FC", x"98FF", x"CD02", x"1106", x"9708", x"7F0A", x"A20B", x"C30B", x"370B", x"9E09", x"3907", x"5604", x"1601", x"25FE", x"B6FB", x"07FA", x"49F9", x"5DF9", x"2AFA", x"62FB", x"A7FC", x"AFFD", x"2DFE", x"03FE", x"42FD", x"00FC", x"A1FA", x"72F9", x"C1F8", x"21F9", x"70FA", x"EAFC", x"5A00", x"DA03", x"6107", x"240A", x"F00B", x"EA0C", x"AA0C", x"910B", x"9209", x"B506", x"A203", x"5B00", x"89FD", x"71FB", x"FCF9", x"92F9", x"BFF9", x"8EFA", x"BAFB", x"C2FC", x"9FFD", x"E3FD", x"7BFD", x"82FC", x"2BFB", x"ACF9", x"71F8", x"A6F7", x"D5F7", x"46F9", x"D2FB", x"D1FF", x"3404", x"7608", x"1B0C", x"330E", x"130F", x"750E", x"680C", x"9E09", x"0C06", x"6702", x"27FF", x"61FC", x"89FA", x"91F9", x"66F9", x"11FA", x"05FB", x"F7FB", x"C4FC", x"EEFC", x"B4FC", x"07FC", x"F7FA", x"CCF9", x"70F8", x"58F7", x"BFF6", x"FAF6", x"A7F8", x"90FB", x"D9FF", x"D604", x"7F09", x"6D0D", x"D00F", x"7F10", x"AB0F", x"6B0D", x"540A", x"F706", x"B703", x"CA00", x"2EFE", x"16FC", x"A5FA", x"05FA", x"FCF9", x"60FA", x"FCFA", x"4AFB", x"38FB", x"FEFA", x"66FA", x"9AFA", x"D6FA", x"7AFB", x"7CFB", x"9CF8", x"F7F6", x"47F7", x"2CFC", x"6902", x"090A", x"0B0E", x"C310", x"EB0F", x"F00C", x"230B", x"2808", x"7E06", x"AF06", x"5404", x"7C03", x"8B03", x"0603", x"D805", x"1801", x"ABFB", x"77ED", x"1CE2", x"00D9", x"2FD4", x"7DD2", x"D7D2", x"2BD3", x"93E0", x"66E4", x"6215", x"9038", x"5D5B", x"EC66", x"2249", x"B429", x"F2EA", x"31D3", x"41BB", x"14D7", x"C8F2", x"271E", x"923B", x"7E3A", x"A224", x"7CFA", x"FBDC", x"83CB", x"27D3", x"C7E2", x"C0F7", x"D9FE", x"9DFE", x"E9E6", x"ABDB", x"B2C6", x"55DF", x"9217", x"873F", x"6F6D", x"F153", x"9D3A", x"FAF2", x"C8CE", x"72B5", x"C7CF", x"2BF4", x"D721", x"E632", x"2230", x"9516", x"B6F3", x"3EDB", x"D9D2", x"5EE2", x"9FF6", x"B406", x"D104", x"A1F7", x"DCE0", x"62CA", x"6DC8", x"A7CB", x"1EF9", x"E839", x"1E56", x"5D6B", x"3535", x"D313", x"14D1", x"12CE", x"FECE", x"5501", x"751B", x"E330", x"231B", x"5DFF", x"7FEA", x"DFE2", x"08EB", x"0BF8", x"6A04", x"A40B", x"0F04", x"20F5", x"78E2", x"A6D6", x"71CF", x"23D4", x"EEE0", x"B8F1", x"D535", x"D341", x"F862", x"6A34", x"881E", x"27E4", x"46DB", x"EDD9", x"20FC", x"7615", x"9422", x"F617", x"F4FB", x"E2F4", x"5DEF", x"10F9", x"70FB", x"F0FF", x"AA00", x"C2FD", x"EDF3", x"41E7", x"61DB", x"E7D1", x"1DD0", x"7ED9", x"20E1", x"3F29", x"C140", x"1D68", x"7443", x"1925", x"6BEA", x"DBD4", x"1AD5", x"F9F3", x"D717", x"8C24", x"7E1E", x"C5FA", x"86F0", x"C1E8", x"04F6", x"38FE", x"C506", x"CE07", x"1302", x"6CF4", x"D4E5", x"D8D7", x"77D3", x"59CE", x"35DE", x"75DB", x"171F", x"8C39", x"725D", x"1F48", x"C626", x"50F8", x"6BD8", x"7EDC", x"FDEF", x"F916", x"AF1D", x"B31D", x"C7F8", x"88EF", x"9AEA", x"76F9", x"3501", x"DE06", x"4805", x"5A00", x"EEF3", x"3DE7", x"F9D9", x"ADD3", x"B9CC", x"BAD7", x"12D6", x"E61B", x"EA3B", x"5463", x"AB4E", x"9A2A", x"BCF9", x"36D6", x"D4DB", x"1CF0", x"D019", x"811F", x"871C", x"10F4", x"96E8", x"D4E5", x"3DFA", x"8407", x"8D0C", x"D209", x"49FF", x"7EF2", x"EEE1", x"D4D9", x"60D1", x"FFCF", x"9BD4", x"05DD", x"FD2A", x"E23E", x"3B69", x"203C", x"5924", x"3DE7", x"CCDC", x"93DC", x"9002", x"D71C", x"6C22", x"FC0D", x"7EEB", x"BDDC", x"A1E7", x"CE04", x"8F17", x"0017", x"5E0A", x"88F7", x"A6E9", x"F2DD", x"27DC", x"CDD6", x"D5DA", x"27D7", x"4FE4", x"8427", x"7238", x"F660", x"4C32", x"8D22", x"E9E4", x"E4E3", x"ABDE", x"EB07", x"5C18", x"8D22", x"BF08", x"7BEB", x"B4D7", x"56E5", x"7507", x"F51B", x"521B", x"3A0A", x"A5F5", x"E4E8", x"08DD", x"36DB", x"D4D5", x"CCD8", x"57CE", x"F9E3", x"2126", x"523C", x"6B64", x"A132", x"A321", x"3FDE", x"E1E2", x"22DD", x"170F", x"4F1D", x"322A", x"F409", x"97E9", x"A8D4", x"E3E2", x"6B02", x"8E1B", x"DD1D", x"CB11", x"3FFB", x"8AED", x"28DF", x"00DD", x"66D4", x"F0D7", x"69CF", x"9AE1", x"FD22", x"5F38", x"E85F", x"B131", x"7C21", x"66E0", x"54E2", x"24DB", x"970A", x"AB1A", x"022A", x"730E", x"F1F2", x"50D7", x"18DF", x"F3FD", x"B817", x"B51E", x"F912", x"3AFF", x"52F0", x"1AE3", x"32DD", x"73D5", x"0AD8", x"C2D0", x"CCDB", x"E81E", x"6733", x"7960", x"A135", x"FB25", x"11E2", x"A5DF", x"91D5", x"C603", x"BA18", x"242D", x"8117", x"5CFA", x"AFDC", x"CDDC", x"73F4", x"D70C", x"A318", x"A416", x"F107", x"62F9", x"7BE5", x"DAD9", x"5FCC", x"F8D0", x"7ACC", x"72E3", x"1425", x"723D", x"EF61", x"3435", x"0321", x"0EE0", x"4ADD", x"F2D4", x"7804", x"6A18", x"E02E", x"5917", x"97FD", x"86DB", x"B6DD", x"31EF", x"EB09", x"8615", x"6C17", x"9F09", x"DAFA", x"15E4", x"09DA", x"11C9", x"00D2", x"06CB", x"12F1", x"0127", x"1943", x"D95B", x"5F32", x"021A", x"CADD", x"07DD", x"7FD7", x"5405", x"EC16", x"B02B", x"2C15", x"0EFE", x"82E3", x"94E5", x"E9F0", x"3F05", x"8B0C", x"CF10", x"B406", x"6BFB", x"72E8", x"8BD9", x"FBCA", x"31CF", x"9BCA", x"030E", x"F427", x"3B59", x"6A46", x"7630", x"E9FB", x"9CDC", x"2CD3", x"43E5", x"BE0A", x"EE20", x"6029", x"C611", x"A5FA", x"14E7", x"A8E6", x"47EF", x"23FE", x"7707", x"0E0E", x"C507", x"5AFA", x"9FE8", x"50D0", x"62CE", x"1FBF", x"F5F5", x"EE1B", x"0C4C", x"1054", x"E03B", x"5C12", x"66E2", x"A5D0", x"53D4", x"4FF9", x"C915", x"EC2C", x"431F", x"A90C", x"FAF1", x"83E7", x"09E5", x"5EEF", x"5EFC", x"1607", x"1F0C", x"E401", x"28F5", x"C2DA", x"14D3", x"A8BB", x"4EEC", x"940E", x"1A44", x"8352", x"7046", x"7D1E", x"8BEE", x"CBD1", x"A0CB", x"9BE9", x"2709", x"AB2A", x"D828", x"361D", x"4000", x"77ED", x"15E1", x"5DE3", x"AEEE", x"4CFE", x"0608", x"2D08", x"F0FA", x"86E6", x"8AD5", x"DCC0", x"9CEB", x"4207", x"7D3F", x"E24A", x"684A", x"1123", x"E6F9", x"52D5", x"42CB", x"73DC", x"30FD", x"891D", x"C42A", x"0628", x"D712", x"ECF9", x"ECE2", x"E7DB", x"D5E0", x"D6F2", x"5C00", x"8B0A", x"D402", x"7EF2", x"26DE", x"91C9", x"C9E9", x"97FD", x"9731", x"563E", x"7F47", x"2829", x"9D09", x"F0E2", x"FFD3", x"52D3", x"5BED", x"8606", x"551F", x"402A", x"B523", x"150C", x"7CF0", x"68DD", x"60D9", x"B7E3", x"D0F3", x"8603", x"FA05", x"A4FF", x"C6E8", x"D3D7", x"D5EA", x"94F7", x"0422", x"CD30", x"7640", x"182E", x"C517", x"9AF4", x"0EE1", x"6BD5", x"3DE2", x"18F5", x"4B11", x"6022", x"6725", x"2615", x"BDFC", x"F7E7", x"A3DD", x"DCDF", x"25EB", x"27FA", x"4703", x"3401", x"58F7", x"65E0", x"4EEC", x"2EF3", x"910F", x"5523", x"B632", x"6D31", x"1D22", x"AC0A", x"3BF3", x"6BE3", x"9DE0", x"DEE8", x"3CFD", x"E20F", x"AE1A", x"E917", x"F809", x"2EF8", x"ECE9", x"48E2", x"4FE5", x"50EE", x"42FB", x"DF00", x"4FFF", x"53F4", x"7EEB", x"7BF4", x"15FC", x"B012", x"D11F", x"D32B", x"D026", x"581C", x"F808", x"59F7", x"AFEA", x"01E8", x"0BEF", x"2AFB", x"6B07", x"F00D", x"F60B", x"C803", x"00F8", x"4CEE", x"A2EA", x"3BED", x"DDF4", x"CCFD", x"E100", x"7C01", x"FCF9", x"9BF0", x"E7F0", x"DEF6", x"1105", x"7F15", x"5120", x"E725", x"2121", x"0F15", x"E905", x"EEF8", x"82F1", x"49EF", x"57F1", x"86F7", x"65FD", x"7601", x"0901", x"D3FC", x"88F8", x"C8F4", x"21F5", x"9AF8", x"DFFC", x"B001", x"7402", x"1400", x"2BFA", x"7FF4", x"71F4", x"16F8", x"5B01", x"D90B", x"1516", x"241A", x"FA1B", x"D016", x"B90F", x"4605", x"EEF9", x"0DF2", x"DFED", x"3BF1", x"DEF7", x"1DFE", x"A901", x"3F00", x"19FD", x"49F8", x"B5F5", x"5BF8", x"2EFA", x"9AFE", x"0900", x"1401", x"AB00", x"9EFE", x"F9FA", x"A0FA", x"F9FB", x"BBFD", x"B203", x"670B", x"BC11", x"1B14", x"580F", x"9907", x"DCFE", x"B4F9", x"1CF9", x"5FFC", x"1F02", x"E304", x"0D05", x"2101", x"11FC", x"F6F7", x"6EF5", x"D2F6", x"2AF9", x"BCFB", x"93FF", x"E801", x"FE01", x"B6FF", x"9BFD", x"66FB", x"CEFA", x"6AFD", x"BC01", x"1E06", x"C506", x"1F03", x"8FFD", x"E8F8", x"8BF7", x"05FA", x"DA00", x"1708", x"9F0A", x"800B", x"8A06", x"3402", x"45FD", x"6AFC", x"61FC", x"35FF", x"D401", x"2504", x"2205", x"4804", x"CC02", x"8800", x"E7FE", x"BAFE", x"9A01", x"3D04", x"5C06", x"CD05", x"E501", x"15FD", x"D8F7", x"FCF5", x"D9F6", x"38FC", x"F100", x"8D03", x"F002", x"2601", x"B5FD", x"43FB", x"57FA", x"5BFB", x"BDFD", x"9D00", x"4D02", x"D803", x"D302", x"1F02", x"7DFF", x"9AFF", x"77FF", x"0B02", x"AC02", x"B904", x"6303", x"8B00", x"A3FD", x"92F8", x"DAF6", x"F6F7", x"D0F9", x"F8FC", x"A8FD", x"9FFD", x"3BFB", x"18FB", x"36FB", x"48FD", x"1200", x"5001", x"7604", x"1B03", x"E202", x"6A01", x"B901", x"7B00", x"3C00", x"2E00", x"3902", x"1006", x"C307", x"4B0A", x"F307", x"A006", x"8604", x"6404", x"7F04", x"F604", x"AF02", x"6801", x"83FB", x"49FA", x"D2F8", x"C0F8", x"ACFB", x"C5FC", x"A2FF", x"41FF", x"3900", x"D4FF", x"9BFF", x"7BFF", x"2A00", x"8301", x"C8FF", x"D600", x"AA00", x"2001", x"5500", x"60FF", x"F8FE", x"9BFC", x"73FD", x"10FD", x"15FE", x"47FE", x"2EFD", x"F7FA", x"3EF9", x"ADF9", x"36FB", x"42FD", x"C2FC", x"B1FE", x"A4FF", x"96FF", x"59FF", x"EFFE", x"2700", x"E700", x"BC01", x"2502", x"E203", x"E602", x"DF05", x"4B06", x"2C06", x"1F07", x"4E07", x"C908", x"D507", x"A70A", x"D607", x"6606", x"A502", x"7FFF", x"9EFE", x"5FFF", x"C9FE", x"FBFC", x"6EFB", x"3EFA", x"8AFA", x"8CFB", x"25FC", x"11FD", x"AEFC", x"D1FA", x"D1FB", x"0CFB", x"9FFC", x"46FD", x"E2FD", x"3EFD", x"0DFD", x"30FE", x"58FE", x"9CFF", x"4800", x"B000", x"9901", x"BBFF", x"F600", x"F901", x"AC02", x"3A03", x"E401", x"1102", x"2400", x"E7FF", x"7700", x"AF01", x"B601", x"8C01", x"1001", x"5901", x"4500", x"A6FF", x"DBFF", x"E5FF", x"2000", x"B200", x"D900", x"1B01", x"2F00", x"AE01", x"FDFF", x"B3FF", x"EDFF", x"62FF", x"CFFF", x"F3FE", x"2201", x"8B00", x"E3FF", x"E0FE", x"C4FE", x"2BFE", x"DDFF", x"AB00", x"5D01", x"2B00", x"72FF", x"73FF", x"18FE", x"21FD", x"F5FD", x"3FFE", x"2CFF", x"E300", x"A7FF", x"9900", x"49FF", x"7EFF", x"D1FF", x"2AFF", x"8F00", x"7F00", x"7D01", x"F700", x"87FF", x"A000", x"BCFF", x"1300", x"CA00", x"3601", x"E601", x"4D02", x"D102", x"7300", x"6DFF", x"20FF", x"A5FE", x"9200", x"6A00", x"2C01", x"9F00", x"D300", x"4DFF", x"84FE", x"E1FD", x"4AFF", x"7AFF", x"0F00", x"C5FF", x"0D01", x"3200", x"9BFF", x"FAFE", x"A4FE", x"44FF", x"09FF", x"7301", x"E900", x"4302", x"D3FF", x"C100", x"5FFE", x"34FE", x"74FE", x"7FFF", x"1A00", x"1300", x"4600", x"CEFF", x"FFFF", x"9100", x"4E00", x"E0FF", x"1900", x"98FF", x"1B00", x"83FF", x"9601", x"E6FF", x"58FF", x"B8FF", x"84FE", x"1700", x"6F00", x"2B01", x"D200", x"9201", x"CEFF", x"B6FE", x"5BFF", x"0300", x"CF00", x"A800", x"2700", x"3600", x"DBFF", x"A300", x"6BFF", x"FAFF", x"8000", x"ECFF", x"6800", x"79FF", x"E100", x"2801", x"A500", x"78FF", x"DDFE", x"B8FE", x"ADFE", x"B4FF", x"C100", x"7D01", x"6601", x"5200", x"EFFE", x"DBFE", x"2CFF", x"1EFF", x"8200", x"42FF", x"EB00", x"B900", x"1000", x"AC00", x"6100", x"2B00", x"52FF", x"FDFF", x"7400", x"8900", x"2E01", x"5A00", x"1600", x"B400", x"A9FF", x"ADFF", x"53FE", x"7BFF", x"3FFF", x"72FF", x"1C00", x"7200", x"1900", x"0400", x"8CFF", x"F8FF", x"71FF", x"ABFF", x"7100", x"FBFF", x"2D00", x"7500", x"82FF", x"DDFF", x"FBFF", x"4D00", x"8F00", x"5000", x"1101", x"C800", x"E6FF", x"7600", x"92FF", x"5500", x"A1FF", x"8D00", x"D5FF", x"2201", x"2DFF", x"BBFF", x"3CFF", x"53FF", x"D1FF", x"A800", x"1200", x"6800", x"DFFF", x"B3FF", x"CCFE", x"EAFF", x"F7FE", x"1100", x"7300", x"5C00", x"E7FF", x"B3FF", x"6000", x"7BFF", x"2300", x"0000", x"BB00", x"7B00", x"A8FF", x"FAFF", x"A3FF", x"9B00", x"3900", x"0001", x"CCFF", x"02FF", x"D3FE", x"DDFF", x"DDFF", x"B800", x"C3FF", x"CF00", x"1300", x"96FF", x"2BFF", x"74FE", x"59FF", x"4900", x"5D01", x"D600", x"4E01", x"3200", x"1F00", x"16FF", x"D6FE", x"59FF", x"0BFF", x"89FF", x"80FF", x"DC00", x"4701", x"DA01", x"9500", x"BFFF", x"1600", x"34FF", x"2600", x"CDFF", x"B800", x"1B00", x"4000", x"F0FE", x"2EFF", x"6AFE", x"54FF", x"5400", x"F700", x"6901", x"D800", x"6800", x"C5FF", x"48FF", x"0100", x"BDFF", x"D6FF", x"2A00", x"DCFF", x"FDFF", x"B7FF", x"C6FF", x"2900", x"B200", x"9800", x"9F00", x"7800", x"1700", x"E7FF", x"DBFF", x"1800", x"0C00", x"82FF", x"7400", x"B0FF", x"C6FF", x"E1FF", x"1400", x"68FF", x"88FF", x"CBFE", x"0400", x"4300", x"9900", x"6900", x"C0FF", x"6BFF", x"BBFF", x"5F00", x"B7FF", x"8A00", x"3000", x"8700", x"1700", x"74FF", x"6FFF", x"2400", x"1A00", x"1000", x"A3FF", x"8C00", x"A9FF", x"5600", x"3E00", x"5300", x"DFFF", x"F7FF", x"73FF", x"FBFF", x"59FF", x"F3FF", x"E0FF", x"B3FF", x"C0FF", x"8400", x"FCFF", x"1101", x"1B00", x"0301", x"C3FF", x"4200", x"BFFF", x"C0FF", x"6FFF", x"7BFF", x"D3FF", x"6000", x"3600", x"D600", x"2A00", x"B5FF", x"B8FF", x"1DFF", x"4D00", x"0D00", x"BC00", x"4300", x"A400", x"7C00", x"A0FF", x"02FF", x"02FF", x"2EFF", x"8AFF", x"D5FF", x"0601", x"CA00", x"9B00", x"0100", x"A4FF", x"2EFF", x"F6FE", x"A9FF", x"F3FF", x"FD00", x"A500", x"9D00", x"8000", x"3B00", x"D5FF", x"3FFF", x"BDFF", x"A7FF", x"DAFF", x"E9FF", x"2B00", x"BA00", x"4400", x"A700", x"46FF", x"A8FF", x"A7FF", x"1900", x"8700", x"5B00", x"5400", x"81FF", x"76FF", x"BFFF", x"F1FF", x"5200", x"A6FF", x"2D00", x"CAFF", x"3600", x"E3FF", x"8800", x"6400", x"4A00", x"D8FF", x"D7FF", x"FFFF", x"CDFF", x"2500", x"66FF", x"E1FF", x"CDFF", x"0000", x"9000", x"0200", x"7200", x"88FF", x"91FF", x"0900", x"3FFF", x"B800", x"E6FF", x"FC00", x"3AFF", x"1600", x"6BFF", x"0A00", x"C2FF", x"62FF", x"7B00", x"7CFF", x"DE00", x"C9FF", x"A700", x"CCFF", x"0800", x"C6FF", x"1900", x"5300", x"9100", x"7200", x"5900", x"E3FF", x"AFFF", x"71FF", x"ADFF", x"1A00", x"6200", x"6B00", x"2C00", x"8FFF", x"4700", x"73FF", x"0C00", x"71FF", x"0700", x"B0FF", x"A400", x"7200", x"3E00", x"FCFF", x"B7FF", x"8FFF", x"46FF", x"D7FF", x"1B00", x"0F01", x"0400", x"D700", x"27FF", x"9FFF", x"08FF", x"0A00", x"7200", x"9B00", x"8F00", x"1900", x"2F00", x"4400", x"9FFF", x"7DFF", x"12FF", x"A1FF", x"0900", x"2400", x"F000", x"AA00", x"9E00", x"F6FE", x"EDFE", x"17FF", x"1100", x"A900", x"3C01", x"1401", x"2900", x"E8FE", x"3FFF", x"3CFF", x"1A00", x"D0FF", x"8300", x"D4FF", x"8D00", x"5200", x"F000", x"7F00", x"2900", x"A7FF", x"E4FE", x"9EFF", x"D9FF", x"F100", x"5200", x"2D00", x"3000", x"D1FF", x"C7FF", x"17FF", x"DBFF", x"E5FF", x"6F00", x"A8FF", x"2E00", x"F7FF", x"3300", x"3700", x"1300", x"D0FF", x"A2FF", x"D9FF", x"4200", x"5D00", x"5400", x"4C00", x"CAFF", x"0E00", x"B4FF", x"DBFF", x"A7FF", x"1400", x"3500", x"5F00", x"3A00", x"4A00", x"1C00", x"44FF", x"19FF", x"D9FE", x"3900", x"9500", x"CA00", x"2600", x"B1FF", x"C7FF", x"B5FF", x"0300", x"C5FF", x"2600", x"E3FF", x"BE00", x"3900", x"B700", x"4F00", x"1300", x"FBFE", x"B5FE", x"10FF", x"3C00", x"F900", x"1001", x"B300", x"1C00", x"B0FF", x"3DFF", x"C5FF", x"FFFF", x"5400", x"7900", x"3300", x"3000", x"9AFF", x"4FFF", x"0AFF", x"BCFF", x"5E00", x"B500", x"6C00", x"1C00", x"EEFF", x"5B00", x"0700", x"B3FF", x"DBFF", x"C5FF", x"FEFF", x"CFFF", x"0D00", x"0200", x"4400", x"F4FF", x"2D00", x"1700", x"1C00", x"5E00", x"3400", x"1600", x"C7FF", x"90FF", x"CAFF", x"EAFF", x"6A00", x"5300", x"2000", x"C2FF", x"79FF", x"D7FF", x"FCFF", x"7200", x"5B00", x"1400", x"B7FF", x"90FF", x"E3FF", x"3600", x"2200", x"1900", x"B6FF", x"EAFF", x"AEFF", x"0300", x"6800", x"5600", x"6900", x"EFFF", x"0400", x"B9FF", x"E7FF", x"C3FF", x"DFFF", x"D0FF", x"F9FF", x"F1FF", x"2600", x"1B00", x"3100", x"F6FF", x"CBFF", x"B5FF", x"D7FF", x"1300", x"4800", x"5800", x"FAFF", x"D2FF", x"B1FF", x"CAFF", x"DDFF", x"E8FF", x"FAFF", x"0200", x"2D00", x"3C00", x"6000", x"5100", x"2A00", x"D2FF", x"AEFF", x"B1FF", x"0700", x"3400", x"3D00", x"2500", x"E6FF", x"E5FF", x"D7FF", x"F5FF", x"1000", x"2200", x"1200", x"DBFF", x"F4FF", x"F7FF", x"4500", x"3800", x"3000", x"F6FF", x"C3FF", x"B4FF", x"D7FF", x"0600", x"2800", x"2F00", x"1600", x"EFFF", x"DCFF", x"EEFF", x"0500", x"1500", x"F5FF", x"0300", x"FAFF", x"0900", x"0500", x"0200", x"0000", x"EFFF", x"F1FF", x"EBFF", x"FFFF", x"1F00", x"3200", x"3300", x"0200", x"E6FF", x"D4FF", x"D3FF", x"E0FF", x"E9FF", x"0B00", x"2200", x"2A00", x"1600", x"F9FF", x"E7FF", x"D6FF", x"EAFF", x"EFFF", x"0800", x"1600", x"2400", x"1600", x"FCFF", x"DFFF", x"E1FF", x"FAFF", x"1600", x"2200", x"2100", x"1400", x"0200", x"EEFF", x"ECFF", x"DFFF", x"DDFF", x"EFFF", x"F5FF", x"0C00", x"0C00", x"0800", x"FEFF", x"0200", x"0C00", x"0E00", x"0D00", x"1000", x"0400", x"0700", x"F9FF", x"FFFF", x"FAFF", x"FFFF", x"FAFF", x"FAFF", x"F9FF", x"0300", x"0700", x"1000", x"0C00", x"1700", x"1A00", x"1400", x"0100", x"EDFF", x"F4FF", x"F1FF", x"F8FF", x"F1FF", x"F2FF", x"F4FF", x"EFFF", x"F0FF", x"FDFF", x"0900", x"1A00", x"1100", x"0900", x"F9FF", x"F3FF", x"F2FF", x"FCFF", x"0200", x"0B00", x"0B00", x"0100", x"FEFF", x"F8FF", x"FAFF", x"F8FF", x"0100", x"0400", x"0600", x"FFFF", x"F6FF", x"F0FF", x"F9FF", x"0100", x"0200", x"0100", x"0100", x"FEFF", x"0300", x"0300", x"0400", x"0200", x"0000", x"0000", x"FBFF", x"FFFF", x"FDFF", x"0200", x"0800", x"0F00", x"1100", x"0D00", x"0700", x"0400", x"0000", x"0000", x"FEFF", x"FFFF", x"FCFF", x"FCFF", x"FCFF", x"0600", x"FEFF", x"FBFF", x"F6FF", x"FDFF", x"FFFF", x"FFFF", x"FFFF", x"0200", x"0700", x"0B00", x"0400", x"FFFF", x"F5FF", x"F7FF", x"F1FF", x"F7FF", x"F7FF", x"FFFF", x"0100", x"0200", x"0200", x"0000", x"0000", x"0200", x"0400", x"0400", x"0700", x"0600", x"0000", x"FBFF", x"F8FF", x"F6FF", x"F5FF", x"F9FF", x"0300", x"0B00", x"1300", x"1100", x"0B00", x"0300", x"FDFF", x"F9FF", x"FDFF", x"0100", x"0400", x"0100", x"FCFF", x"FAFF", x"F7FF", x"F8FF", x"F8FF", x"F9FF", x"FBFF", x"0000", x"0400", x"0700", x"0600", x"0300", x"0000", x"FDFF", x"0100", x"0100", x"0200", x"0300", x"0400", x"0100", x"0100", x"0000", x"FCFF", x"FBFF", x"FAFF", x"FAFF", x"FBFF", x"FFFF", x"0300", x"0500", x"0200", x"0000", x"FEFF", x"0100", x"0300", x"0500", x"0200", x"FEFF", x"0000", x"FDFF", x"0100", x"FFFF", x"0300", x"0200", x"0100", x"FDFF", x"FCFF", x"FFFF", x"0200", x"0400", x"0300", x"0300", x"0300", x"0300", x"0500", x"0700", x"0500", x"0200", x"0000", x"FEFF", x"FAFF", x"FCFF", x"FDFF", x"0100", x"0200", x"0300", x"FFFF", x"FEFF", x"0100", x"0000", x"FFFF", x"FEFF", x"FCFF", x"FCFF", x"FEFF", x"0100", x"FFFF", x"FEFF", x"FEFF", x"FCFF", x"FAFF", x"F8FF", x"FCFF", x"FDFF", x"0000", x"FFFF", x"0100", x"0200", x"0300", x"0200", x"0200", x"0400", x"0300", x"0500", x"0400", x"0200", x"FFFF", x"FEFF", x"0000", x"0000", x"0000", x"0000", x"0100", x"0000", x"0100", x"0200", x"0400", x"0600", x"0500", x"0400", x"0100", x"FBFF", x"FCFF", x"FBFF", x"FEFF", x"FEFF", x"FFFF", x"0000", x"FFFF", x"FDFF", x"FDFF", x"0100", x"0400", x"0700", x"0700", x"0500", x"0200", x"FFFF", x"FEFF", x"FDFF", x"FDFF", x"FEFF", x"0000", x"0000", x"0000", x"FFFF", x"FEFF", x"0000", x"0000", x"FEFF", x"FEFF", x"FFFF", x"FFFF", x"0000", x"0000", x"0100", x"0000", x"0000", x"FEFF", x"FDFF", x"FBFF", x"FCFF", x"FEFF", x"0000", x"0100", x"FFFF", x"FBFF", x"FDFF", x"FEFF", x"FEFF", x"0000", x"FFFF", x"FFFF", x"0200", x"0200", x"0200", x"0100", x"0100", x"0100", x"0100", x"0300", x"0300", x"0000", x"0200", x"0200", x"0200", x"0000", x"0200", x"0300", x"0200", x"0300", x"0200", x"0100", x"0100", x"FEFF", x"FFFF", x"FDFF", x"FEFF", x"0000", x"FDFF", x"FFFF", x"FEFF", x"FFFF", x"FEFF", x"FEFF", x"0000", x"0100", x"0200", x"0200", x"0000", x"0000", x"0000", x"0000", x"0200", x"0200", x"0100", x"0100", x"0000", x"FFFF", x"FFFF", x"0000", x"FEFF", x"0000", x"0200", x"0200", x"0300", x"0200", x"0200", x"0200", x"0100", x"0100", x"0100", x"0100", x"0200", x"0300", x"0100", x"0100", x"0000", x"FFFF", x"0000", x"0000", x"FFFF", x"0000", x"0000", x"0100", x"0000", x"FEFF", x"FFFF", x"FFFF", x"0100", x"0300", x"0300", x"0200", x"0000", x"0100", x"FFFF", x"FEFF", x"FFFF", x"FDFF", x"FDFF", x"FEFF", x"FEFF", x"FEFF", x"FFFF", x"FDFF", x"FCFF", x"FDFF", x"FEFF", x"0000", x"0000", x"0100", x"0000", x"0000", x"0000", x"0000", x"0100", x"0000", x"FFFF", x"FFFF", x"0000", x"FFFF", x"0000", x"0000", x"0000", x"0100", x"0300", x"0600", x"0600", x"0600", x"0400", x"0300", x"0100", x"0100", x"0000", x"FFFF", x"FCFF", x"FCFF", x"FBFF", x"FAFF", x"FAFF", x"FCFF", x"FDFF", x"FCFF", x"FCFF", x"FEFF", x"FFFF", x"0000", x"0000", x"0100", x"0200", x"0000", x"0100", x"0200", x"0300", x"0200", x"0200", x"0100", x"FEFF", x"FEFF", x"FFFF", x"FFFF", x"0100", x"0000", x"0100", x"0000", x"FFFF", x"0000", x"0200", x"0200", x"0200", x"0200", x"0200", x"0200", x"0200", x"0200", x"0200", x"0100", x"0100", x"0100", x"0100", x"0300", x"0200", x"0200", x"0200", x"0200", x"0300", x"0200", x"0300", x"0300", x"0200", x"0000", x"0100", x"0000", x"FFFF", x"FEFF", x"FFFF", x"FFFF", x"FEFF", x"FFFF", x"FEFF", x"FEFF", x"FEFF", x"FEFF", x"FDFF", x"FCFF", x"FCFF", x"FDFF", x"FDFF", x"FFFF", x"FFFF", x"FEFF", x"FDFF", x"FFFF", x"0000", x"0100", x"FEFF", x"FFFF", x"FCFF", x"0200", x"0300", x"FCFF", x"F9FF", x"FCFF", x"0300", x"0200", x"0100", x"0300", x"0800", x"0600", x"0200", x"0100", x"0100", x"0100", x"FFFF", x"FAFF", x"F7FF", x"F7FF", x"F7FF", x"F7FF", x"F8FF", x"F9FF", x"FBFF", x"FEFF", x"FEFF", x"FFFF", x"0000", x"0200", x"0200", x"0300", x"0400", x"0500", x"0500", x"0400", x"0400", x"0400", x"0500", x"0600", x"0700", x"0600", x"0600", x"0800", x"0800", x"0900", x"0900", x"0900", x"0800", x"0900", x"0800", x"0700", x"0400", x"0100", x"0200", x"0100", x"0200", x"0000", x"0000", x"0100", x"0200", x"0100", x"FFFF", x"FCFF", x"FCFF", x"F9FF", x"F8FF", x"F9FF", x"FAFF", x"FAFF", x"FAFF", x"FAFF", x"F9FF", x"F9FF", x"F8FF", x"F8FF", x"F8FF", x"F8FF", x"FAFF", x"F9FF", x"FAFF", x"FCFF", x"FCFF", x"FBFF", x"FAFF", x"FBFF", x"FCFF", x"FCFF", x"FDFF", x"FDFF", x"FCFF", x"FCFF", x"FBFF", x"FCFF", x"FDFF", x"0000", x"0100", x"0300", x"0400", x"0300", x"0400", x"0400", x"0200", x"0200", x"0400", x"0400", x"0300", x"0200", x"0200", x"0300", x"0300", x"0300", x"0400", x"0400", x"0400", x"0600", x"0600", x"0800", x"0900", x"0900", x"0700", x"0400", x"0300", x"0100", x"0200", x"0300", x"0400", x"0400", x"0400", x"0400", x"0300", x"0400", x"0200", x"0400", x"0500", x"0400", x"0400", x"0100", x"0100", x"0100", x"FFFF", x"FEFF", x"FCFF", x"FDFF", x"FDFF", x"FDFF", x"FEFF", x"FEFF", x"FDFF", x"FDFF", x"FEFF", x"0000", x"0100", x"0000", x"0000", x"0100", x"0000", x"FFFF", x"FFFF", x"FFFF", x"FCFF", x"FEFF", x"FCFF", x"FCFF", x"FDFF", x"FDFF", x"FDFF", x"FEFF", x"FBFF", x"FBFF", x"FAFF", x"FBFF", x"FBFF", x"FAFF", x"FAFF", x"FBFF", x"FBFF", x"F9FF", x"FAFF", x"FAFF", x"FCFF", x"FEFF", x"FFFF", x"0000", x"FFFF", x"0100", x"0000", x"FFFF", x"0000", x"0000", x"FFFF", x"0000", x"FFFF", x"0000", x"0000", x"0100", x"0300", x"0300", x"0100", x"0200", x"0400", x"0400", x"0600", x"0500", x"0500", x"0500", x"0500", x"0500", x"0500", x"0500", x"0500");
				--
				
				signal DATA		  : STD_LOGIC_VECTOR (15 downto 0);
			--	signal DATA1	  : STD_LOGIC_VECTOR (15 downto 0);
				signal DATA2	  : STD_LOGIC_VECTOR (15 downto 0);
				signal BIG_DATA  : STD_LOGIC_VECTOR (15 downto 0);
				signal DAC_DATA  : STD_LOGIC_VECTOR (15 downto 0);
				signal DAC_REG   : STD_LOGIC_VECTOR (31 downto 0);
				signal SEND		  : STD_LOGIC  :='1';
				signal SENDING   : STD_LOGIC  :='0';
				signal SCK_CLK	  : STD_LOGIC  ;
				signal FF_ONE    : STD_LOGIC  :='0';
			--	signal FF_ZERO   : STD_LOGIC  :='0';
				signal FF_BES    : STD_LOGIC  :='0';
				signal DIVCNTR   : integer    :=0;
				signal SDATA     : integer;
				signal UDATA     : integer;
				signal i         : integer range 0 to 5403:=0;
			--	signal k         : integer range 0 to 4846:=0;
				signal j         : integer range 0 to 4660:=0;
begin
				
		DAC_CLR<='1';
		FPGA_INIT_B<='1';
		SF_CE0<='1';
		AD_CONV<='0';
		AMP_CS<='1';
		SPI_SS_B<='1';
		
		CLKDIV:  process(CLK) is begin											 
					 if(rising_edge(CLK)) then										
						if(DIVCNTR>=391) then DIVCNTR <=0; SCK_CLK<='1'; 		
						else DIVCNTR <= DIVCNTR +1; SCK_CLK<='0';  end if;
					 end if;
					end process;	
				
			DAC:	process(SCK_CLK) is
						variable COUNTER : integer range 0 to 31 := 0;	
					begin
			
				if rising_edge(SCK_CLK) then
					if(B_ONE='1') then FF_ONE<='1'; FF_BES<='0'; 
					--elsif(B_ZERO='1') then FF_ZERO<='1'; FF_ONE<='0'; 
					elsif(B_BES='1') then FF_BES<='1'; FF_ONE<='0'; end if; 
					
					DATA <=One_voice(i);
				 --DATA1<=Zero_voice(k);
					DATA2<=Bes_voice(j);
					
					if(SEND = '1') then
						if(FF_ONE='1') then	
							BIG_DATA <= DATA(7 downto 0) & DATA(15 downto 8);
							SDATA <= conv_integer(signed(BIG_DATA));
							UDATA <= SDATA + 32768;
							DAC_DATA <= CONV_STD_LOGIC_VECTOR(UDATA,16);
							DAC_REG <=  "00000000" & "0011" & "1111" & DAC_DATA(15 downto 4) & "0000" ;
							COUNTER := 0;	
							DAC_CS <= '0';
							SENDING <= '1';
							SEND <= '0';
							i<=i+1; 
--						elsif(FF_ZERO='1') then
--							BIG_DATA <= DATA1(7 downto 0) & DATA1(15 downto 8);
--							SDATA <= conv_integer(signed(BIG_DATA));
--							UDATA <= SDATA + 32768;
--							DAC_DATA <= CONV_STD_LOGIC_VECTOR(UDATA,16);
--							DAC_REG <=  "00000000" & "0011" & "1111" & DAC_DATA(15 downto 4) & "0000" ;
--							COUNTER := 0;	
--							DAC_CS <= '0';
--							SENDING <= '1';
--							SEND <= '0';
--							k<=k+1; 
						elsif(FF_BES='1') then
							BIG_DATA <= DATA2(7 downto 0) & DATA2(15 downto 8);
							SDATA <= conv_integer(signed(BIG_DATA));
							UDATA <= SDATA + 32768;
							DAC_DATA <= CONV_STD_LOGIC_VECTOR(UDATA,16);
							DAC_REG <=  "00000000" & "0011" & "1111" & DAC_DATA(15 downto 4) & "0000" ;
							COUNTER := 0;	
							DAC_CS <= '0';
							SENDING <= '1';
							SEND <= '0';
							j<=j+1; end if;	
						end if;
					
						if SENDING = '1' then	
							DAC_REG(31 downto 1) <= DAC_REG(30 downto 0); 
										
								if (COUNTER = 31) then		
									COUNTER := 0;	
									DAC_CS <= '1';
									SENDING <= '0'; 
									SEND <= '1';
								else
									COUNTER := COUNTER + 1;	
								end if;
						end if;	
						
							
				end if;
						
				end process;
				SPI_MOSI <= DAC_REG(31);
				SPI_SCK  <= SCK_CLK;
end Behavioral;

